/**
 *  @file   bch_45_32.vh
 *  @brief  (27,16)BCH符号
 *
 *  @par    Copyright
 *  (C) 2012 Taichi Ishitani All Rights Reserved.
 *
 *  @author Taichi Ishitani
 *
 *  @date   0.0.00  2012/05/01  T. Ishitani     coding start
 */

function [12:0] f_calc_parity_bch_45_32 (
    input   [31:0]  i_d
);
    f_calc_parity_bch_45_32 = {
        //  x^31 +   x^30 +   x^29 +   x^28 +   x^27 +   x^26 +   x^25 +   x^24 +   x^23 +   x^22 +   x^21 +   x^20 +   x^19 +   x^18 +   x^17 +   x^16 +   x^15 +   x^14 +   x^13 +   x^12 +   x^11 +   x^10 +   x^9 +   x^8 +   x^7 +   x^6 +   x^5 +   x^4 +   x^3 +   x^2 +   x^1 +   x^0
        ^{                  i_d[29], i_d[28],          i_d[26], i_d[25], i_d[24], i_d[23], i_d[22], i_d[21],                   i_d[18],                   i_d[15],                   i_d[12], i_d[11], i_d[10],         i_d[8],         i_d[6], i_d[5],                         i_d[1]        },    // 0x37e49d62
        ^{                           i_d[28], i_d[27],          i_d[25], i_d[24], i_d[23], i_d[22], i_d[21], i_d[20],                   i_d[17],                   i_d[14],                   i_d[11], i_d[10], i_d[9],         i_d[7],         i_d[5], i_d[4],                         i_d[0]},    // 0x1bf24eb1
        ^{i_d[31],          i_d[29], i_d[28], i_d[27],          i_d[25],                                     i_d[20], i_d[19], i_d[18],          i_d[16], i_d[15],          i_d[13], i_d[12], i_d[11],          i_d[9],                         i_d[5], i_d[4], i_d[3],         i_d[1]        },    // 0xba1dba3a
        ^{i_d[31], i_d[30],          i_d[28], i_d[27], i_d[26],          i_d[24],                                     i_d[19], i_d[18], i_d[17],          i_d[15], i_d[14],          i_d[12], i_d[11], i_d[10],         i_d[8],                         i_d[4], i_d[3], i_d[2],         i_d[0]},    // 0xdd0edd1d
        ^{i_d[31], i_d[30],          i_d[28], i_d[27],                   i_d[24],          i_d[22], i_d[21],                            i_d[17], i_d[16], i_d[15], i_d[14], i_d[13], i_d[12],                   i_d[9], i_d[8], i_d[7], i_d[6], i_d[5],         i_d[3], i_d[2]                },    // 0xd963f3ec
        ^{i_d[31], i_d[30], i_d[29],          i_d[27], i_d[26],                   i_d[23],          i_d[21], i_d[20],                            i_d[16], i_d[15], i_d[14], i_d[13], i_d[12], i_d[11],                  i_d[8], i_d[7], i_d[6], i_d[5], i_d[4], i_d[2],         i_d[1]        },    // 0xecb1f9f6
        ^{i_d[31], i_d[30], i_d[29], i_d[28],          i_d[26], i_d[25],                   i_d[22],          i_d[20], i_d[19],                            i_d[15], i_d[14], i_d[13], i_d[12], i_d[11], i_d[10],                 i_d[7], i_d[6], i_d[5], i_d[4], i_d[3],         i_d[1], i_d[0]},    // 0xf658fcfb
        ^{         i_d[30],                   i_d[27], i_d[26],                   i_d[23], i_d[22],                   i_d[19],                            i_d[15], i_d[14], i_d[13],                            i_d[9], i_d[8],                         i_d[4], i_d[3], i_d[2], i_d[1], i_d[0]},    // 0x4cc8e31f
        ^{                           i_d[28],                            i_d[24], i_d[23],                                                                i_d[15], i_d[14], i_d[13],          i_d[11], i_d[10],                 i_d[7], i_d[6], i_d[5],         i_d[3], i_d[2],         i_d[0]},    // 0x1180eced
        ^{i_d[31],          i_d[29], i_d[28], i_d[27], i_d[26], i_d[25], i_d[24],                   i_d[21],                   i_d[18],                   i_d[15], i_d[14], i_d[13],          i_d[11],          i_d[9], i_d[8],                         i_d[4],         i_d[2]                },    // 0xbf24eb14
        ^{i_d[31], i_d[30],          i_d[28], i_d[27], i_d[26], i_d[25], i_d[24], i_d[23],                   i_d[20],                   i_d[17],                   i_d[14], i_d[13], i_d[12],          i_d[10],         i_d[8], i_d[7],                         i_d[3],         i_d[1]        },    // 0xdf92758a
        ^{         i_d[30], i_d[29],          i_d[27], i_d[26], i_d[25], i_d[24], i_d[23], i_d[22],                   i_d[19],                   i_d[16],                   i_d[13], i_d[12], i_d[11],          i_d[9],         i_d[7], i_d[6],                         i_d[2],         i_d[0]},    // 0x6fc93ac5
        ^{                  i_d[29],                   i_d[26],          i_d[24],          i_d[22],                            i_d[18], i_d[17], i_d[16],                            i_d[12],          i_d[10], i_d[9],                 i_d[6],                                 i_d[1], i_d[0]}     // 0x25471643
    };
endfunction

function [1034:0] f_decode_syndrome_bch_45_32 (
    input   [12:0]  i_syn
);
    f_decode_syndrome_bch_45_32 = {
        ((i_syn == 13'h042a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1307) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1890) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0862) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1523) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b82) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1cd3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1f7a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1eaf) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1e44) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b08) ? 1'b1 : 1'b0),
        ((i_syn == 13'h01ae) ? 1'b1 : 1'b0),
        ((i_syn == 13'h11c5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0cc9) ? 1'b1 : 1'b0),
        ((i_syn == 13'h024f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1034) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0c30) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0232) ? 1'b1 : 1'b0),
        ((i_syn == 13'h100b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1916) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d99) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ae7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1460) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0e1a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h161f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1a1c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0924) ? 1'b1 : 1'b0),
        ((i_syn == 13'h00b8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0476) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1329) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0dbf) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17cc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0fcc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03cc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h05cc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h06cc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h074c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h078c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h07ec) ? 1'b1 : 1'b0),
        ((i_syn == 13'h07dc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h07c4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h07c8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h07ce) ? 1'b1 : 1'b0),
        ((i_syn == 13'h07cd) ? 1'b1 : 1'b0),
        ((i_syn == 13'h172d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1cba) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0c48) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1109) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1fa8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h18f9) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b50) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1a85) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1a6e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0f22) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0584) ? 1'b1 : 1'b0),
        ((i_syn == 13'h15ef) ? 1'b1 : 1'b0),
        ((i_syn == 13'h08e3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0665) ? 1'b1 : 1'b0),
        ((i_syn == 13'h141e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h081a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0618) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1421) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d3c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h19b3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ecd) ? 1'b1 : 1'b0),
        ((i_syn == 13'h104a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a30) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1235) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1e36) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d0e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0492) ? 1'b1 : 1'b0),
        ((i_syn == 13'h005c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1703) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0995) ? 1'b1 : 1'b0),
        ((i_syn == 13'h13e6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0be6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h07e6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h01e6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h02e6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0366) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03a6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03c6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03f6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03ee) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03e2) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03e4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03e7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b97) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b65) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0624) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0885) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0fd4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0c7d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0da8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d43) ? 1'b1 : 1'b0),
        ((i_syn == 13'h180f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h12a9) ? 1'b1 : 1'b0),
        ((i_syn == 13'h02c2) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1fce) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1148) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0333) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1f37) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1135) ? 1'b1 : 1'b0),
        ((i_syn == 13'h030c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a11) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0e9e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h19e0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0767) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d1d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0518) ? 1'b1 : 1'b0),
        ((i_syn == 13'h091b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1a23) ? 1'b1 : 1'b0),
        ((i_syn == 13'h13bf) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1771) ? 1'b1 : 1'b0),
        ((i_syn == 13'h002e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1eb8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h04cb) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1ccb) ? 1'b1 : 1'b0),
        ((i_syn == 13'h10cb) ? 1'b1 : 1'b0),
        ((i_syn == 13'h16cb) ? 1'b1 : 1'b0),
        ((i_syn == 13'h15cb) ? 1'b1 : 1'b0),
        ((i_syn == 13'h144b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h148b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14eb) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14db) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14c3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14cf) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14c9) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14ca) ? 1'b1 : 1'b0),
        ((i_syn == 13'h10f2) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0db3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0312) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0443) ? 1'b1 : 1'b0),
        ((i_syn == 13'h07ea) ? 1'b1 : 1'b0),
        ((i_syn == 13'h063f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h06d4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1398) ? 1'b1 : 1'b0),
        ((i_syn == 13'h193e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0955) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1459) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1adf) ? 1'b1 : 1'b0),
        ((i_syn == 13'h08a4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14a0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1aa2) ? 1'b1 : 1'b0),
        ((i_syn == 13'h089b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0186) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0509) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1277) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0cf0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h168a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0e8f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h028c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h11b4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1828) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1ce6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0bb9) ? 1'b1 : 1'b0),
        ((i_syn == 13'h152f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0f5c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h175c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b5c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d5c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1e5c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1fdc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1f1c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1f7c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1f4c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1f54) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1f58) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1f5e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1f5d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d41) ? 1'b1 : 1'b0),
        ((i_syn == 13'h13e0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14b1) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1718) ? 1'b1 : 1'b0),
        ((i_syn == 13'h16cd) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1626) ? 1'b1 : 1'b0),
        ((i_syn == 13'h036a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h09cc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h19a7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h04ab) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a2d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1856) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0452) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a50) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1869) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1174) ? 1'b1 : 1'b0),
        ((i_syn == 13'h15fb) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0285) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1c02) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0678) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1e7d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h127e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0146) ? 1'b1 : 1'b0),
        ((i_syn == 13'h08da) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0c14) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b4b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h05dd) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1fae) ? 1'b1 : 1'b0),
        ((i_syn == 13'h07ae) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0bae) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0dae) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0eae) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0f2e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0fee) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0f8e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0fbe) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0fa6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0faa) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0fac) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0faf) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ea1) ? 1'b1 : 1'b0),
        ((i_syn == 13'h09f0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a59) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b8c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b67) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1e2b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h148d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h04e6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h19ea) ? 1'b1 : 1'b0),
        ((i_syn == 13'h176c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0517) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1913) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1711) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0528) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0c35) ? 1'b1 : 1'b0),
        ((i_syn == 13'h08ba) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1fc4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0143) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b39) ? 1'b1 : 1'b0),
        ((i_syn == 13'h033c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0f3f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1c07) ? 1'b1 : 1'b0),
        ((i_syn == 13'h159b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1155) ? 1'b1 : 1'b0),
        ((i_syn == 13'h060a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h189c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h02ef) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1aef) ? 1'b1 : 1'b0),
        ((i_syn == 13'h16ef) ? 1'b1 : 1'b0),
        ((i_syn == 13'h10ef) ? 1'b1 : 1'b0),
        ((i_syn == 13'h13ef) ? 1'b1 : 1'b0),
        ((i_syn == 13'h126f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h12af) ? 1'b1 : 1'b0),
        ((i_syn == 13'h12cf) ? 1'b1 : 1'b0),
        ((i_syn == 13'h12ff) ? 1'b1 : 1'b0),
        ((i_syn == 13'h12e7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h12eb) ? 1'b1 : 1'b0),
        ((i_syn == 13'h12ed) ? 1'b1 : 1'b0),
        ((i_syn == 13'h12ee) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0751) ? 1'b1 : 1'b0),
        ((i_syn == 13'h04f8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h052d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h05c6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h108a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1a2c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a47) ? 1'b1 : 1'b0),
        ((i_syn == 13'h174b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h19cd) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0bb6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17b2) ? 1'b1 : 1'b0),
        ((i_syn == 13'h19b0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b89) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0294) ? 1'b1 : 1'b0),
        ((i_syn == 13'h061b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1165) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0fe2) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1598) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d9d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h019e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h12a6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b3a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1ff4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h08ab) ? 1'b1 : 1'b0),
        ((i_syn == 13'h163d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0c4e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h144e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h184e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1e4e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d4e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1cce) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1c0e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1c6e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1c5e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1c46) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1c4a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1c4c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1c4f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03a9) ? 1'b1 : 1'b0),
        ((i_syn == 13'h027c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0297) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17db) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d7d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d16) ? 1'b1 : 1'b0),
        ((i_syn == 13'h101a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1e9c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ce7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h10e3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1ee1) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0cd8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h05c5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h014a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1634) ? 1'b1 : 1'b0),
        ((i_syn == 13'h08b3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h12c9) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0acc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h06cf) ? 1'b1 : 1'b0),
        ((i_syn == 13'h15f7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1c6b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h18a5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ffa) ? 1'b1 : 1'b0),
        ((i_syn == 13'h116c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b1f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h131f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1f1f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h191f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1a1f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b9f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b5f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b3f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b0f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b17) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b1b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b1d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b1e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h01d5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h013e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1472) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1ed4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ebf) ? 1'b1 : 1'b0),
        ((i_syn == 13'h13b3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d35) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0f4e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h134a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d48) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0f71) ? 1'b1 : 1'b0),
        ((i_syn == 13'h066c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h02e3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h159d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b1a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1160) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0965) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0566) ? 1'b1 : 1'b0),
        ((i_syn == 13'h165e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1fc2) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b0c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0c53) ? 1'b1 : 1'b0),
        ((i_syn == 13'h12c5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h08b6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h10b6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1cb6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1ab6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h19b6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1836) ? 1'b1 : 1'b0),
        ((i_syn == 13'h18f6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1896) ? 1'b1 : 1'b0),
        ((i_syn == 13'h18a6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h18be) ? 1'b1 : 1'b0),
        ((i_syn == 13'h18b2) ? 1'b1 : 1'b0),
        ((i_syn == 13'h18b4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h18b7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h00eb) ? 1'b1 : 1'b0),
        ((i_syn == 13'h15a7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1f01) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0f6a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1266) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1ce0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0e9b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h129f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1c9d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ea4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h07b9) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0336) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1448) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0acf) ? 1'b1 : 1'b0),
        ((i_syn == 13'h10b5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h08b0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h04b3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h178b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1e17) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1ad9) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d86) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1310) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0963) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1163) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d63) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b63) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1863) ? 1'b1 : 1'b0),
        ((i_syn == 13'h19e3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1923) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1943) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1973) ? 1'b1 : 1'b0),
        ((i_syn == 13'h196b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1967) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1961) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1962) ? 1'b1 : 1'b0),
        ((i_syn == 13'h154c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1fea) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0f81) ? 1'b1 : 1'b0),
        ((i_syn == 13'h128d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1c0b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0e70) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1274) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1c76) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0e4f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0752) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03dd) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14a3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a24) ? 1'b1 : 1'b0),
        ((i_syn == 13'h105e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h085b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0458) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1760) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1efc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1a32) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d6d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h13fb) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0988) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1188) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d88) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b88) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1888) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1908) ? 1'b1 : 1'b0),
        ((i_syn == 13'h19c8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h19a8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1998) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1980) ? 1'b1 : 1'b0),
        ((i_syn == 13'h198c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h198a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1989) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0aa6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1acd) ? 1'b1 : 1'b0),
        ((i_syn == 13'h07c1) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0947) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b3c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0738) ? 1'b1 : 1'b0),
        ((i_syn == 13'h093a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b03) ? 1'b1 : 1'b0),
        ((i_syn == 13'h121e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1691) ? 1'b1 : 1'b0),
        ((i_syn == 13'h01ef) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1f68) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0512) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d17) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1114) ? 1'b1 : 1'b0),
        ((i_syn == 13'h022c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0bb0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0f7e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1821) ? 1'b1 : 1'b0),
        ((i_syn == 13'h06b7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1cc4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h04c4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h08c4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ec4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0dc4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0c44) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0c84) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ce4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0cd4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ccc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0cc0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0cc6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0cc5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h106b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d67) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03e1) ? 1'b1 : 1'b0),
        ((i_syn == 13'h119a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d9e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h039c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h11a5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h18b8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1c37) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b49) ? 1'b1 : 1'b0),
        ((i_syn == 13'h15ce) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0fb4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17b1) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1bb2) ? 1'b1 : 1'b0),
        ((i_syn == 13'h088a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0116) ? 1'b1 : 1'b0),
        ((i_syn == 13'h05d8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1287) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0c11) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1662) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0e62) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0262) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0462) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0762) ? 1'b1 : 1'b0),
        ((i_syn == 13'h06e2) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0622) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0642) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0672) ? 1'b1 : 1'b0),
        ((i_syn == 13'h066a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0666) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0660) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0663) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d0c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h138a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h01f1) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1df5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h13f7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h01ce) ? 1'b1 : 1'b0),
        ((i_syn == 13'h08d3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0c5c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b22) ? 1'b1 : 1'b0),
        ((i_syn == 13'h05a5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1fdf) ? 1'b1 : 1'b0),
        ((i_syn == 13'h07da) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0bd9) ? 1'b1 : 1'b0),
        ((i_syn == 13'h18e1) ? 1'b1 : 1'b0),
        ((i_syn == 13'h117d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h15b3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h02ec) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1c7a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0609) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1e09) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1209) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1409) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1709) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1689) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1649) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1629) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1619) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1601) ? 1'b1 : 1'b0),
        ((i_syn == 13'h160d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h160b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1608) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0e86) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1cfd) ? 1'b1 : 1'b0),
        ((i_syn == 13'h00f9) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0efb) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1cc2) ? 1'b1 : 1'b0),
        ((i_syn == 13'h15df) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1150) ? 1'b1 : 1'b0),
        ((i_syn == 13'h062e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h18a9) ? 1'b1 : 1'b0),
        ((i_syn == 13'h02d3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1ad6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h16d5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h05ed) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0c71) ? 1'b1 : 1'b0),
        ((i_syn == 13'h08bf) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1fe0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0176) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b05) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0305) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0f05) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0905) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a05) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b85) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b45) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b25) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b15) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b0d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b01) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b07) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b04) ? 1'b1 : 1'b0),
        ((i_syn == 13'h127b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0e7f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h007d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1244) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b59) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1fd6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h08a8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h162f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0c55) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1450) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1853) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b6b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h02f7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0639) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1166) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ff0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1583) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d83) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0183) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0783) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0483) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0503) ? 1'b1 : 1'b0),
        ((i_syn == 13'h05c3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h05a3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0593) ? 1'b1 : 1'b0),
        ((i_syn == 13'h058b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0587) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0581) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0582) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1c04) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1206) ? 1'b1 : 1'b0),
        ((i_syn == 13'h003f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0922) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0dad) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1ad3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0454) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1e2e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h062b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a28) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1910) ? 1'b1 : 1'b0),
        ((i_syn == 13'h108c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1442) ? 1'b1 : 1'b0),
        ((i_syn == 13'h031d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d8b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h07f8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1ff8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h13f8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h15f8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h16f8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1778) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17b8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17d8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17e8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17f0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17fc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17fa) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17f9) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0e02) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1c3b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1526) ? 1'b1 : 1'b0),
        ((i_syn == 13'h11a9) ? 1'b1 : 1'b0),
        ((i_syn == 13'h06d7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1850) ? 1'b1 : 1'b0),
        ((i_syn == 13'h022a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1a2f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h162c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0514) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0c88) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0846) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1f19) ? 1'b1 : 1'b0),
        ((i_syn == 13'h018f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1bfc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03fc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ffc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h09fc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0afc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b7c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0bbc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0bdc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0bec) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0bf4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0bf8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0bfe) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0bfd) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1239) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b24) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1fab) ? 1'b1 : 1'b0),
        ((i_syn == 13'h08d5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1652) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0c28) ? 1'b1 : 1'b0),
        ((i_syn == 13'h142d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h182e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b16) ? 1'b1 : 1'b0),
        ((i_syn == 13'h028a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0644) ? 1'b1 : 1'b0),
        ((i_syn == 13'h111b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0f8d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h15fe) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0dfe) ? 1'b1 : 1'b0),
        ((i_syn == 13'h01fe) ? 1'b1 : 1'b0),
        ((i_syn == 13'h07fe) ? 1'b1 : 1'b0),
        ((i_syn == 13'h04fe) ? 1'b1 : 1'b0),
        ((i_syn == 13'h057e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h05be) ? 1'b1 : 1'b0),
        ((i_syn == 13'h05de) ? 1'b1 : 1'b0),
        ((i_syn == 13'h05ee) ? 1'b1 : 1'b0),
        ((i_syn == 13'h05f6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h05fa) ? 1'b1 : 1'b0),
        ((i_syn == 13'h05fc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h05ff) ? 1'b1 : 1'b0),
        ((i_syn == 13'h091d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d92) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1aec) ? 1'b1 : 1'b0),
        ((i_syn == 13'h046b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1e11) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0614) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a17) ? 1'b1 : 1'b0),
        ((i_syn == 13'h192f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h10b3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h147d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0322) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1db4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h07c7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1fc7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h13c7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h15c7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h16c7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1747) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1787) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17e7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17d7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17cf) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17c3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17c5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17c6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h048f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h13f1) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d76) ? 1'b1 : 1'b0),
        ((i_syn == 13'h170c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0f09) ? 1'b1 : 1'b0),
        ((i_syn == 13'h030a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1032) ? 1'b1 : 1'b0),
        ((i_syn == 13'h19ae) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d60) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a3f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14a9) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0eda) ? 1'b1 : 1'b0),
        ((i_syn == 13'h16da) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1ada) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1cda) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1fda) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1e5a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1e9a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1efa) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1eca) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1ed2) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1ede) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1ed8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1edb) ? 1'b1 : 1'b0),
        ((i_syn == 13'h177e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h09f9) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1383) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b86) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0785) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14bd) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d21) ? 1'b1 : 1'b0),
        ((i_syn == 13'h19ef) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0eb0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1026) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a55) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1255) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1e55) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1855) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b55) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1ad5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1a15) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1a75) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1a45) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1a5d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1a51) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1a57) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1a54) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1e87) ? 1'b1 : 1'b0),
        ((i_syn == 13'h04fd) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1cf8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h10fb) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03c3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a5f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0e91) ? 1'b1 : 1'b0),
        ((i_syn == 13'h19ce) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0758) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d2b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h052b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h092b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0f2b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0c2b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0dab) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d6b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d0b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d3b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d23) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d2f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d29) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d2a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1a7a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h027f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0e7c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d44) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14d8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1016) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0749) ? 1'b1 : 1'b0),
        ((i_syn == 13'h19df) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03ac) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1bac) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17ac) ? 1'b1 : 1'b0),
        ((i_syn == 13'h11ac) ? 1'b1 : 1'b0),
        ((i_syn == 13'h12ac) ? 1'b1 : 1'b0),
        ((i_syn == 13'h132c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h13ec) ? 1'b1 : 1'b0),
        ((i_syn == 13'h138c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h13bc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h13a4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h13a8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h13ae) ? 1'b1 : 1'b0),
        ((i_syn == 13'h13ad) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1805) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1406) ? 1'b1 : 1'b0),
        ((i_syn == 13'h073e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ea2) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a6c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d33) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03a5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h19d6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h01d6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0dd6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0bd6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h08d6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0956) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0996) ? 1'b1 : 1'b0),
        ((i_syn == 13'h09f6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h09c6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h09de) ? 1'b1 : 1'b0),
        ((i_syn == 13'h09d2) ? 1'b1 : 1'b0),
        ((i_syn == 13'h09d4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h09d7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0c03) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1f3b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h16a7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1269) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0536) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1ba0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h01d3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h19d3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h15d3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h13d3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h10d3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1153) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1193) ? 1'b1 : 1'b0),
        ((i_syn == 13'h11f3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h11c3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h11db) ? 1'b1 : 1'b0),
        ((i_syn == 13'h11d7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h11d1) ? 1'b1 : 1'b0),
        ((i_syn == 13'h11d2) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1338) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1aa4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1e6a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0935) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17a3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0dd0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h15d0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h19d0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1fd0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1cd0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d50) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1d90) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1df0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1dc0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1dd8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1dd4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1dd2) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1dd1) ? 1'b1 : 1'b0),
        ((i_syn == 13'h099c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d52) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1a0d) ? 1'b1 : 1'b0),
        ((i_syn == 13'h049b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1ee8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h06e8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ae8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ce8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0fe8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0e68) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ea8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ec8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ef8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ee0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0eec) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0eea) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ee9) ? 1'b1 : 1'b0),
        ((i_syn == 13'h04ce) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1391) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d07) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1774) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0f74) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0374) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0574) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0674) ? 1'b1 : 1'b0),
        ((i_syn == 13'h07f4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0734) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0754) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0764) ? 1'b1 : 1'b0),
        ((i_syn == 13'h077c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0770) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0776) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0775) ? 1'b1 : 1'b0),
        ((i_syn == 13'h175f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h09c9) ? 1'b1 : 1'b0),
        ((i_syn == 13'h13ba) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0bba) ? 1'b1 : 1'b0),
        ((i_syn == 13'h07ba) ? 1'b1 : 1'b0),
        ((i_syn == 13'h01ba) ? 1'b1 : 1'b0),
        ((i_syn == 13'h02ba) ? 1'b1 : 1'b0),
        ((i_syn == 13'h033a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03fa) ? 1'b1 : 1'b0),
        ((i_syn == 13'h039a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03aa) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03b2) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03be) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03b8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03bb) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1e96) ? 1'b1 : 1'b0),
        ((i_syn == 13'h04e5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1ce5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h10e5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h16e5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h15e5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1465) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14a5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14c5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14f5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14ed) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14e1) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14e7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14e4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1a73) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0273) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0e73) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0873) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b73) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0af3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a33) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a53) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a63) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a7b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a77) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a71) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a72) ? 1'b1 : 1'b0),
        ((i_syn == 13'h07cc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03e6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14cb) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1f5c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0fae) ? 1'b1 : 1'b0),
        ((i_syn == 13'h12ef) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1c4e) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1b1f) ? 1'b1 : 1'b0),
        ((i_syn == 13'h18b6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1963) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1988) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0cc4) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0662) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1609) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0b05) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0583) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17f8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0bfc) ? 1'b1 : 1'b0),
        ((i_syn == 13'h05fe) ? 1'b1 : 1'b0),
        ((i_syn == 13'h17c7) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1eda) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1a55) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0d2b) ? 1'b1 : 1'b0),
        ((i_syn == 13'h13ac) ? 1'b1 : 1'b0),
        ((i_syn == 13'h09d6) ? 1'b1 : 1'b0),
        ((i_syn == 13'h11d3) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1dd0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0ee8) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0774) ? 1'b1 : 1'b0),
        ((i_syn == 13'h03ba) ? 1'b1 : 1'b0),
        ((i_syn == 13'h14e5) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a73) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1800) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1400) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1200) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1100) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1080) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1040) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1020) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1010) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1008) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1004) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1002) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1001) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0c00) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0a00) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0900) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0880) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0840) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0820) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0810) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0808) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0804) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0802) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0801) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0600) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0500) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0480) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0440) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0420) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0410) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0408) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0404) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0402) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0401) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0300) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0280) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0240) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0220) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0210) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0208) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0204) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0202) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0201) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0180) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0140) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0120) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0110) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0108) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0104) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0102) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0101) ? 1'b1 : 1'b0),
        ((i_syn == 13'h00c0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h00a0) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0090) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0088) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0084) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0082) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0081) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0060) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0050) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0048) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0044) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0042) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0041) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0030) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0028) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0024) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0022) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0021) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0018) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0014) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0012) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0011) ? 1'b1 : 1'b0),
        ((i_syn == 13'h000c) ? 1'b1 : 1'b0),
        ((i_syn == 13'h000a) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0009) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0006) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0005) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0003) ? 1'b1 : 1'b0),
        ((i_syn == 13'h1000) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0800) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0400) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0200) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0100) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0080) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0040) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0020) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0010) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0008) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0004) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0002) ? 1'b1 : 1'b0),
        ((i_syn == 13'h0001) ? 1'b1 : 1'b0)
    };
endfunction

function [31:0] f_select_pattern_bch_45_32 (
    input   [943:0] i_sel
);
    f_select_pattern_bch_45_32  = ({32{i_sel[943]}} & 32'hc0000000)     //  syndrome : 0x042a
                                | ({32{i_sel[942]}} & 32'ha0000000)     //  syndrome : 0x1307
                                | ({32{i_sel[941]}} & 32'h90000000)     //  syndrome : 0x1890
                                | ({32{i_sel[940]}} & 32'h88000000)     //  syndrome : 0x0862
                                | ({32{i_sel[939]}} & 32'h84000000)     //  syndrome : 0x1523
                                | ({32{i_sel[938]}} & 32'h82000000)     //  syndrome : 0x1b82
                                | ({32{i_sel[937]}} & 32'h81000000)     //  syndrome : 0x1cd3
                                | ({32{i_sel[936]}} & 32'h80800000)     //  syndrome : 0x1f7a
                                | ({32{i_sel[935]}} & 32'h80400000)     //  syndrome : 0x1eaf
                                | ({32{i_sel[934]}} & 32'h80200000)     //  syndrome : 0x1e44
                                | ({32{i_sel[933]}} & 32'h80100000)     //  syndrome : 0x0b08
                                | ({32{i_sel[932]}} & 32'h80080000)     //  syndrome : 0x01ae
                                | ({32{i_sel[931]}} & 32'h80040000)     //  syndrome : 0x11c5
                                | ({32{i_sel[930]}} & 32'h80020000)     //  syndrome : 0x0cc9
                                | ({32{i_sel[929]}} & 32'h80010000)     //  syndrome : 0x024f
                                | ({32{i_sel[928]}} & 32'h80008000)     //  syndrome : 0x1034
                                | ({32{i_sel[927]}} & 32'h80004000)     //  syndrome : 0x0c30
                                | ({32{i_sel[926]}} & 32'h80002000)     //  syndrome : 0x0232
                                | ({32{i_sel[925]}} & 32'h80001000)     //  syndrome : 0x100b
                                | ({32{i_sel[924]}} & 32'h80000800)     //  syndrome : 0x1916
                                | ({32{i_sel[923]}} & 32'h80000400)     //  syndrome : 0x1d99
                                | ({32{i_sel[922]}} & 32'h80000200)     //  syndrome : 0x0ae7
                                | ({32{i_sel[921]}} & 32'h80000100)     //  syndrome : 0x1460
                                | ({32{i_sel[920]}} & 32'h80000080)     //  syndrome : 0x0e1a
                                | ({32{i_sel[919]}} & 32'h80000040)     //  syndrome : 0x161f
                                | ({32{i_sel[918]}} & 32'h80000020)     //  syndrome : 0x1a1c
                                | ({32{i_sel[917]}} & 32'h80000010)     //  syndrome : 0x0924
                                | ({32{i_sel[916]}} & 32'h80000008)     //  syndrome : 0x00b8
                                | ({32{i_sel[915]}} & 32'h80000004)     //  syndrome : 0x0476
                                | ({32{i_sel[914]}} & 32'h80000002)     //  syndrome : 0x1329
                                | ({32{i_sel[913]}} & 32'h80000001)     //  syndrome : 0x0dbf
                                | ({32{i_sel[912]}} & 32'h80000000)     //  syndrome : 0x17cc
                                | ({32{i_sel[911]}} & 32'h80000000)     //  syndrome : 0x0fcc
                                | ({32{i_sel[910]}} & 32'h80000000)     //  syndrome : 0x03cc
                                | ({32{i_sel[909]}} & 32'h80000000)     //  syndrome : 0x05cc
                                | ({32{i_sel[908]}} & 32'h80000000)     //  syndrome : 0x06cc
                                | ({32{i_sel[907]}} & 32'h80000000)     //  syndrome : 0x074c
                                | ({32{i_sel[906]}} & 32'h80000000)     //  syndrome : 0x078c
                                | ({32{i_sel[905]}} & 32'h80000000)     //  syndrome : 0x07ec
                                | ({32{i_sel[904]}} & 32'h80000000)     //  syndrome : 0x07dc
                                | ({32{i_sel[903]}} & 32'h80000000)     //  syndrome : 0x07c4
                                | ({32{i_sel[902]}} & 32'h80000000)     //  syndrome : 0x07c8
                                | ({32{i_sel[901]}} & 32'h80000000)     //  syndrome : 0x07ce
                                | ({32{i_sel[900]}} & 32'h80000000)     //  syndrome : 0x07cd
                                | ({32{i_sel[899]}} & 32'h60000000)     //  syndrome : 0x172d
                                | ({32{i_sel[898]}} & 32'h50000000)     //  syndrome : 0x1cba
                                | ({32{i_sel[897]}} & 32'h48000000)     //  syndrome : 0x0c48
                                | ({32{i_sel[896]}} & 32'h44000000)     //  syndrome : 0x1109
                                | ({32{i_sel[895]}} & 32'h42000000)     //  syndrome : 0x1fa8
                                | ({32{i_sel[894]}} & 32'h41000000)     //  syndrome : 0x18f9
                                | ({32{i_sel[893]}} & 32'h40800000)     //  syndrome : 0x1b50
                                | ({32{i_sel[892]}} & 32'h40400000)     //  syndrome : 0x1a85
                                | ({32{i_sel[891]}} & 32'h40200000)     //  syndrome : 0x1a6e
                                | ({32{i_sel[890]}} & 32'h40100000)     //  syndrome : 0x0f22
                                | ({32{i_sel[889]}} & 32'h40080000)     //  syndrome : 0x0584
                                | ({32{i_sel[888]}} & 32'h40040000)     //  syndrome : 0x15ef
                                | ({32{i_sel[887]}} & 32'h40020000)     //  syndrome : 0x08e3
                                | ({32{i_sel[886]}} & 32'h40010000)     //  syndrome : 0x0665
                                | ({32{i_sel[885]}} & 32'h40008000)     //  syndrome : 0x141e
                                | ({32{i_sel[884]}} & 32'h40004000)     //  syndrome : 0x081a
                                | ({32{i_sel[883]}} & 32'h40002000)     //  syndrome : 0x0618
                                | ({32{i_sel[882]}} & 32'h40001000)     //  syndrome : 0x1421
                                | ({32{i_sel[881]}} & 32'h40000800)     //  syndrome : 0x1d3c
                                | ({32{i_sel[880]}} & 32'h40000400)     //  syndrome : 0x19b3
                                | ({32{i_sel[879]}} & 32'h40000200)     //  syndrome : 0x0ecd
                                | ({32{i_sel[878]}} & 32'h40000100)     //  syndrome : 0x104a
                                | ({32{i_sel[877]}} & 32'h40000080)     //  syndrome : 0x0a30
                                | ({32{i_sel[876]}} & 32'h40000040)     //  syndrome : 0x1235
                                | ({32{i_sel[875]}} & 32'h40000020)     //  syndrome : 0x1e36
                                | ({32{i_sel[874]}} & 32'h40000010)     //  syndrome : 0x0d0e
                                | ({32{i_sel[873]}} & 32'h40000008)     //  syndrome : 0x0492
                                | ({32{i_sel[872]}} & 32'h40000004)     //  syndrome : 0x005c
                                | ({32{i_sel[871]}} & 32'h40000002)     //  syndrome : 0x1703
                                | ({32{i_sel[870]}} & 32'h40000001)     //  syndrome : 0x0995
                                | ({32{i_sel[869]}} & 32'h40000000)     //  syndrome : 0x13e6
                                | ({32{i_sel[868]}} & 32'h40000000)     //  syndrome : 0x0be6
                                | ({32{i_sel[867]}} & 32'h40000000)     //  syndrome : 0x07e6
                                | ({32{i_sel[866]}} & 32'h40000000)     //  syndrome : 0x01e6
                                | ({32{i_sel[865]}} & 32'h40000000)     //  syndrome : 0x02e6
                                | ({32{i_sel[864]}} & 32'h40000000)     //  syndrome : 0x0366
                                | ({32{i_sel[863]}} & 32'h40000000)     //  syndrome : 0x03a6
                                | ({32{i_sel[862]}} & 32'h40000000)     //  syndrome : 0x03c6
                                | ({32{i_sel[861]}} & 32'h40000000)     //  syndrome : 0x03f6
                                | ({32{i_sel[860]}} & 32'h40000000)     //  syndrome : 0x03ee
                                | ({32{i_sel[859]}} & 32'h40000000)     //  syndrome : 0x03e2
                                | ({32{i_sel[858]}} & 32'h40000000)     //  syndrome : 0x03e4
                                | ({32{i_sel[857]}} & 32'h40000000)     //  syndrome : 0x03e7
                                | ({32{i_sel[856]}} & 32'h30000000)     //  syndrome : 0x0b97
                                | ({32{i_sel[855]}} & 32'h28000000)     //  syndrome : 0x1b65
                                | ({32{i_sel[854]}} & 32'h24000000)     //  syndrome : 0x0624
                                | ({32{i_sel[853]}} & 32'h22000000)     //  syndrome : 0x0885
                                | ({32{i_sel[852]}} & 32'h21000000)     //  syndrome : 0x0fd4
                                | ({32{i_sel[851]}} & 32'h20800000)     //  syndrome : 0x0c7d
                                | ({32{i_sel[850]}} & 32'h20400000)     //  syndrome : 0x0da8
                                | ({32{i_sel[849]}} & 32'h20200000)     //  syndrome : 0x0d43
                                | ({32{i_sel[848]}} & 32'h20100000)     //  syndrome : 0x180f
                                | ({32{i_sel[847]}} & 32'h20080000)     //  syndrome : 0x12a9
                                | ({32{i_sel[846]}} & 32'h20040000)     //  syndrome : 0x02c2
                                | ({32{i_sel[845]}} & 32'h20020000)     //  syndrome : 0x1fce
                                | ({32{i_sel[844]}} & 32'h20010000)     //  syndrome : 0x1148
                                | ({32{i_sel[843]}} & 32'h20008000)     //  syndrome : 0x0333
                                | ({32{i_sel[842]}} & 32'h20004000)     //  syndrome : 0x1f37
                                | ({32{i_sel[841]}} & 32'h20002000)     //  syndrome : 0x1135
                                | ({32{i_sel[840]}} & 32'h20001000)     //  syndrome : 0x030c
                                | ({32{i_sel[839]}} & 32'h20000800)     //  syndrome : 0x0a11
                                | ({32{i_sel[838]}} & 32'h20000400)     //  syndrome : 0x0e9e
                                | ({32{i_sel[837]}} & 32'h20000200)     //  syndrome : 0x19e0
                                | ({32{i_sel[836]}} & 32'h20000100)     //  syndrome : 0x0767
                                | ({32{i_sel[835]}} & 32'h20000080)     //  syndrome : 0x1d1d
                                | ({32{i_sel[834]}} & 32'h20000040)     //  syndrome : 0x0518
                                | ({32{i_sel[833]}} & 32'h20000020)     //  syndrome : 0x091b
                                | ({32{i_sel[832]}} & 32'h20000010)     //  syndrome : 0x1a23
                                | ({32{i_sel[831]}} & 32'h20000008)     //  syndrome : 0x13bf
                                | ({32{i_sel[830]}} & 32'h20000004)     //  syndrome : 0x1771
                                | ({32{i_sel[829]}} & 32'h20000002)     //  syndrome : 0x002e
                                | ({32{i_sel[828]}} & 32'h20000001)     //  syndrome : 0x1eb8
                                | ({32{i_sel[827]}} & 32'h20000000)     //  syndrome : 0x04cb
                                | ({32{i_sel[826]}} & 32'h20000000)     //  syndrome : 0x1ccb
                                | ({32{i_sel[825]}} & 32'h20000000)     //  syndrome : 0x10cb
                                | ({32{i_sel[824]}} & 32'h20000000)     //  syndrome : 0x16cb
                                | ({32{i_sel[823]}} & 32'h20000000)     //  syndrome : 0x15cb
                                | ({32{i_sel[822]}} & 32'h20000000)     //  syndrome : 0x144b
                                | ({32{i_sel[821]}} & 32'h20000000)     //  syndrome : 0x148b
                                | ({32{i_sel[820]}} & 32'h20000000)     //  syndrome : 0x14eb
                                | ({32{i_sel[819]}} & 32'h20000000)     //  syndrome : 0x14db
                                | ({32{i_sel[818]}} & 32'h20000000)     //  syndrome : 0x14c3
                                | ({32{i_sel[817]}} & 32'h20000000)     //  syndrome : 0x14cf
                                | ({32{i_sel[816]}} & 32'h20000000)     //  syndrome : 0x14c9
                                | ({32{i_sel[815]}} & 32'h20000000)     //  syndrome : 0x14ca
                                | ({32{i_sel[814]}} & 32'h18000000)     //  syndrome : 0x10f2
                                | ({32{i_sel[813]}} & 32'h14000000)     //  syndrome : 0x0db3
                                | ({32{i_sel[812]}} & 32'h12000000)     //  syndrome : 0x0312
                                | ({32{i_sel[811]}} & 32'h11000000)     //  syndrome : 0x0443
                                | ({32{i_sel[810]}} & 32'h10800000)     //  syndrome : 0x07ea
                                | ({32{i_sel[809]}} & 32'h10400000)     //  syndrome : 0x063f
                                | ({32{i_sel[808]}} & 32'h10200000)     //  syndrome : 0x06d4
                                | ({32{i_sel[807]}} & 32'h10100000)     //  syndrome : 0x1398
                                | ({32{i_sel[806]}} & 32'h10080000)     //  syndrome : 0x193e
                                | ({32{i_sel[805]}} & 32'h10040000)     //  syndrome : 0x0955
                                | ({32{i_sel[804]}} & 32'h10020000)     //  syndrome : 0x1459
                                | ({32{i_sel[803]}} & 32'h10010000)     //  syndrome : 0x1adf
                                | ({32{i_sel[802]}} & 32'h10008000)     //  syndrome : 0x08a4
                                | ({32{i_sel[801]}} & 32'h10004000)     //  syndrome : 0x14a0
                                | ({32{i_sel[800]}} & 32'h10002000)     //  syndrome : 0x1aa2
                                | ({32{i_sel[799]}} & 32'h10001000)     //  syndrome : 0x089b
                                | ({32{i_sel[798]}} & 32'h10000800)     //  syndrome : 0x0186
                                | ({32{i_sel[797]}} & 32'h10000400)     //  syndrome : 0x0509
                                | ({32{i_sel[796]}} & 32'h10000200)     //  syndrome : 0x1277
                                | ({32{i_sel[795]}} & 32'h10000100)     //  syndrome : 0x0cf0
                                | ({32{i_sel[794]}} & 32'h10000080)     //  syndrome : 0x168a
                                | ({32{i_sel[793]}} & 32'h10000040)     //  syndrome : 0x0e8f
                                | ({32{i_sel[792]}} & 32'h10000020)     //  syndrome : 0x028c
                                | ({32{i_sel[791]}} & 32'h10000010)     //  syndrome : 0x11b4
                                | ({32{i_sel[790]}} & 32'h10000008)     //  syndrome : 0x1828
                                | ({32{i_sel[789]}} & 32'h10000004)     //  syndrome : 0x1ce6
                                | ({32{i_sel[788]}} & 32'h10000002)     //  syndrome : 0x0bb9
                                | ({32{i_sel[787]}} & 32'h10000001)     //  syndrome : 0x152f
                                | ({32{i_sel[786]}} & 32'h10000000)     //  syndrome : 0x0f5c
                                | ({32{i_sel[785]}} & 32'h10000000)     //  syndrome : 0x175c
                                | ({32{i_sel[784]}} & 32'h10000000)     //  syndrome : 0x1b5c
                                | ({32{i_sel[783]}} & 32'h10000000)     //  syndrome : 0x1d5c
                                | ({32{i_sel[782]}} & 32'h10000000)     //  syndrome : 0x1e5c
                                | ({32{i_sel[781]}} & 32'h10000000)     //  syndrome : 0x1fdc
                                | ({32{i_sel[780]}} & 32'h10000000)     //  syndrome : 0x1f1c
                                | ({32{i_sel[779]}} & 32'h10000000)     //  syndrome : 0x1f7c
                                | ({32{i_sel[778]}} & 32'h10000000)     //  syndrome : 0x1f4c
                                | ({32{i_sel[777]}} & 32'h10000000)     //  syndrome : 0x1f54
                                | ({32{i_sel[776]}} & 32'h10000000)     //  syndrome : 0x1f58
                                | ({32{i_sel[775]}} & 32'h10000000)     //  syndrome : 0x1f5e
                                | ({32{i_sel[774]}} & 32'h10000000)     //  syndrome : 0x1f5d
                                | ({32{i_sel[773]}} & 32'h0c000000)     //  syndrome : 0x1d41
                                | ({32{i_sel[772]}} & 32'h0a000000)     //  syndrome : 0x13e0
                                | ({32{i_sel[771]}} & 32'h09000000)     //  syndrome : 0x14b1
                                | ({32{i_sel[770]}} & 32'h08800000)     //  syndrome : 0x1718
                                | ({32{i_sel[769]}} & 32'h08400000)     //  syndrome : 0x16cd
                                | ({32{i_sel[768]}} & 32'h08200000)     //  syndrome : 0x1626
                                | ({32{i_sel[767]}} & 32'h08100000)     //  syndrome : 0x036a
                                | ({32{i_sel[766]}} & 32'h08080000)     //  syndrome : 0x09cc
                                | ({32{i_sel[765]}} & 32'h08040000)     //  syndrome : 0x19a7
                                | ({32{i_sel[764]}} & 32'h08020000)     //  syndrome : 0x04ab
                                | ({32{i_sel[763]}} & 32'h08010000)     //  syndrome : 0x0a2d
                                | ({32{i_sel[762]}} & 32'h08008000)     //  syndrome : 0x1856
                                | ({32{i_sel[761]}} & 32'h08004000)     //  syndrome : 0x0452
                                | ({32{i_sel[760]}} & 32'h08002000)     //  syndrome : 0x0a50
                                | ({32{i_sel[759]}} & 32'h08001000)     //  syndrome : 0x1869
                                | ({32{i_sel[758]}} & 32'h08000800)     //  syndrome : 0x1174
                                | ({32{i_sel[757]}} & 32'h08000400)     //  syndrome : 0x15fb
                                | ({32{i_sel[756]}} & 32'h08000200)     //  syndrome : 0x0285
                                | ({32{i_sel[755]}} & 32'h08000100)     //  syndrome : 0x1c02
                                | ({32{i_sel[754]}} & 32'h08000080)     //  syndrome : 0x0678
                                | ({32{i_sel[753]}} & 32'h08000040)     //  syndrome : 0x1e7d
                                | ({32{i_sel[752]}} & 32'h08000020)     //  syndrome : 0x127e
                                | ({32{i_sel[751]}} & 32'h08000010)     //  syndrome : 0x0146
                                | ({32{i_sel[750]}} & 32'h08000008)     //  syndrome : 0x08da
                                | ({32{i_sel[749]}} & 32'h08000004)     //  syndrome : 0x0c14
                                | ({32{i_sel[748]}} & 32'h08000002)     //  syndrome : 0x1b4b
                                | ({32{i_sel[747]}} & 32'h08000001)     //  syndrome : 0x05dd
                                | ({32{i_sel[746]}} & 32'h08000000)     //  syndrome : 0x1fae
                                | ({32{i_sel[745]}} & 32'h08000000)     //  syndrome : 0x07ae
                                | ({32{i_sel[744]}} & 32'h08000000)     //  syndrome : 0x0bae
                                | ({32{i_sel[743]}} & 32'h08000000)     //  syndrome : 0x0dae
                                | ({32{i_sel[742]}} & 32'h08000000)     //  syndrome : 0x0eae
                                | ({32{i_sel[741]}} & 32'h08000000)     //  syndrome : 0x0f2e
                                | ({32{i_sel[740]}} & 32'h08000000)     //  syndrome : 0x0fee
                                | ({32{i_sel[739]}} & 32'h08000000)     //  syndrome : 0x0f8e
                                | ({32{i_sel[738]}} & 32'h08000000)     //  syndrome : 0x0fbe
                                | ({32{i_sel[737]}} & 32'h08000000)     //  syndrome : 0x0fa6
                                | ({32{i_sel[736]}} & 32'h08000000)     //  syndrome : 0x0faa
                                | ({32{i_sel[735]}} & 32'h08000000)     //  syndrome : 0x0fac
                                | ({32{i_sel[734]}} & 32'h08000000)     //  syndrome : 0x0faf
                                | ({32{i_sel[733]}} & 32'h06000000)     //  syndrome : 0x0ea1
                                | ({32{i_sel[732]}} & 32'h05000000)     //  syndrome : 0x09f0
                                | ({32{i_sel[731]}} & 32'h04800000)     //  syndrome : 0x0a59
                                | ({32{i_sel[730]}} & 32'h04400000)     //  syndrome : 0x0b8c
                                | ({32{i_sel[729]}} & 32'h04200000)     //  syndrome : 0x0b67
                                | ({32{i_sel[728]}} & 32'h04100000)     //  syndrome : 0x1e2b
                                | ({32{i_sel[727]}} & 32'h04080000)     //  syndrome : 0x148d
                                | ({32{i_sel[726]}} & 32'h04040000)     //  syndrome : 0x04e6
                                | ({32{i_sel[725]}} & 32'h04020000)     //  syndrome : 0x19ea
                                | ({32{i_sel[724]}} & 32'h04010000)     //  syndrome : 0x176c
                                | ({32{i_sel[723]}} & 32'h04008000)     //  syndrome : 0x0517
                                | ({32{i_sel[722]}} & 32'h04004000)     //  syndrome : 0x1913
                                | ({32{i_sel[721]}} & 32'h04002000)     //  syndrome : 0x1711
                                | ({32{i_sel[720]}} & 32'h04001000)     //  syndrome : 0x0528
                                | ({32{i_sel[719]}} & 32'h04000800)     //  syndrome : 0x0c35
                                | ({32{i_sel[718]}} & 32'h04000400)     //  syndrome : 0x08ba
                                | ({32{i_sel[717]}} & 32'h04000200)     //  syndrome : 0x1fc4
                                | ({32{i_sel[716]}} & 32'h04000100)     //  syndrome : 0x0143
                                | ({32{i_sel[715]}} & 32'h04000080)     //  syndrome : 0x1b39
                                | ({32{i_sel[714]}} & 32'h04000040)     //  syndrome : 0x033c
                                | ({32{i_sel[713]}} & 32'h04000020)     //  syndrome : 0x0f3f
                                | ({32{i_sel[712]}} & 32'h04000010)     //  syndrome : 0x1c07
                                | ({32{i_sel[711]}} & 32'h04000008)     //  syndrome : 0x159b
                                | ({32{i_sel[710]}} & 32'h04000004)     //  syndrome : 0x1155
                                | ({32{i_sel[709]}} & 32'h04000002)     //  syndrome : 0x060a
                                | ({32{i_sel[708]}} & 32'h04000001)     //  syndrome : 0x189c
                                | ({32{i_sel[707]}} & 32'h04000000)     //  syndrome : 0x02ef
                                | ({32{i_sel[706]}} & 32'h04000000)     //  syndrome : 0x1aef
                                | ({32{i_sel[705]}} & 32'h04000000)     //  syndrome : 0x16ef
                                | ({32{i_sel[704]}} & 32'h04000000)     //  syndrome : 0x10ef
                                | ({32{i_sel[703]}} & 32'h04000000)     //  syndrome : 0x13ef
                                | ({32{i_sel[702]}} & 32'h04000000)     //  syndrome : 0x126f
                                | ({32{i_sel[701]}} & 32'h04000000)     //  syndrome : 0x12af
                                | ({32{i_sel[700]}} & 32'h04000000)     //  syndrome : 0x12cf
                                | ({32{i_sel[699]}} & 32'h04000000)     //  syndrome : 0x12ff
                                | ({32{i_sel[698]}} & 32'h04000000)     //  syndrome : 0x12e7
                                | ({32{i_sel[697]}} & 32'h04000000)     //  syndrome : 0x12eb
                                | ({32{i_sel[696]}} & 32'h04000000)     //  syndrome : 0x12ed
                                | ({32{i_sel[695]}} & 32'h04000000)     //  syndrome : 0x12ee
                                | ({32{i_sel[694]}} & 32'h03000000)     //  syndrome : 0x0751
                                | ({32{i_sel[693]}} & 32'h02800000)     //  syndrome : 0x04f8
                                | ({32{i_sel[692]}} & 32'h02400000)     //  syndrome : 0x052d
                                | ({32{i_sel[691]}} & 32'h02200000)     //  syndrome : 0x05c6
                                | ({32{i_sel[690]}} & 32'h02100000)     //  syndrome : 0x108a
                                | ({32{i_sel[689]}} & 32'h02080000)     //  syndrome : 0x1a2c
                                | ({32{i_sel[688]}} & 32'h02040000)     //  syndrome : 0x0a47
                                | ({32{i_sel[687]}} & 32'h02020000)     //  syndrome : 0x174b
                                | ({32{i_sel[686]}} & 32'h02010000)     //  syndrome : 0x19cd
                                | ({32{i_sel[685]}} & 32'h02008000)     //  syndrome : 0x0bb6
                                | ({32{i_sel[684]}} & 32'h02004000)     //  syndrome : 0x17b2
                                | ({32{i_sel[683]}} & 32'h02002000)     //  syndrome : 0x19b0
                                | ({32{i_sel[682]}} & 32'h02001000)     //  syndrome : 0x0b89
                                | ({32{i_sel[681]}} & 32'h02000800)     //  syndrome : 0x0294
                                | ({32{i_sel[680]}} & 32'h02000400)     //  syndrome : 0x061b
                                | ({32{i_sel[679]}} & 32'h02000200)     //  syndrome : 0x1165
                                | ({32{i_sel[678]}} & 32'h02000100)     //  syndrome : 0x0fe2
                                | ({32{i_sel[677]}} & 32'h02000080)     //  syndrome : 0x1598
                                | ({32{i_sel[676]}} & 32'h02000040)     //  syndrome : 0x0d9d
                                | ({32{i_sel[675]}} & 32'h02000020)     //  syndrome : 0x019e
                                | ({32{i_sel[674]}} & 32'h02000010)     //  syndrome : 0x12a6
                                | ({32{i_sel[673]}} & 32'h02000008)     //  syndrome : 0x1b3a
                                | ({32{i_sel[672]}} & 32'h02000004)     //  syndrome : 0x1ff4
                                | ({32{i_sel[671]}} & 32'h02000002)     //  syndrome : 0x08ab
                                | ({32{i_sel[670]}} & 32'h02000001)     //  syndrome : 0x163d
                                | ({32{i_sel[669]}} & 32'h02000000)     //  syndrome : 0x0c4e
                                | ({32{i_sel[668]}} & 32'h02000000)     //  syndrome : 0x144e
                                | ({32{i_sel[667]}} & 32'h02000000)     //  syndrome : 0x184e
                                | ({32{i_sel[666]}} & 32'h02000000)     //  syndrome : 0x1e4e
                                | ({32{i_sel[665]}} & 32'h02000000)     //  syndrome : 0x1d4e
                                | ({32{i_sel[664]}} & 32'h02000000)     //  syndrome : 0x1cce
                                | ({32{i_sel[663]}} & 32'h02000000)     //  syndrome : 0x1c0e
                                | ({32{i_sel[662]}} & 32'h02000000)     //  syndrome : 0x1c6e
                                | ({32{i_sel[661]}} & 32'h02000000)     //  syndrome : 0x1c5e
                                | ({32{i_sel[660]}} & 32'h02000000)     //  syndrome : 0x1c46
                                | ({32{i_sel[659]}} & 32'h02000000)     //  syndrome : 0x1c4a
                                | ({32{i_sel[658]}} & 32'h02000000)     //  syndrome : 0x1c4c
                                | ({32{i_sel[657]}} & 32'h02000000)     //  syndrome : 0x1c4f
                                | ({32{i_sel[656]}} & 32'h01800000)     //  syndrome : 0x03a9
                                | ({32{i_sel[655]}} & 32'h01400000)     //  syndrome : 0x027c
                                | ({32{i_sel[654]}} & 32'h01200000)     //  syndrome : 0x0297
                                | ({32{i_sel[653]}} & 32'h01100000)     //  syndrome : 0x17db
                                | ({32{i_sel[652]}} & 32'h01080000)     //  syndrome : 0x1d7d
                                | ({32{i_sel[651]}} & 32'h01040000)     //  syndrome : 0x0d16
                                | ({32{i_sel[650]}} & 32'h01020000)     //  syndrome : 0x101a
                                | ({32{i_sel[649]}} & 32'h01010000)     //  syndrome : 0x1e9c
                                | ({32{i_sel[648]}} & 32'h01008000)     //  syndrome : 0x0ce7
                                | ({32{i_sel[647]}} & 32'h01004000)     //  syndrome : 0x10e3
                                | ({32{i_sel[646]}} & 32'h01002000)     //  syndrome : 0x1ee1
                                | ({32{i_sel[645]}} & 32'h01001000)     //  syndrome : 0x0cd8
                                | ({32{i_sel[644]}} & 32'h01000800)     //  syndrome : 0x05c5
                                | ({32{i_sel[643]}} & 32'h01000400)     //  syndrome : 0x014a
                                | ({32{i_sel[642]}} & 32'h01000200)     //  syndrome : 0x1634
                                | ({32{i_sel[641]}} & 32'h01000100)     //  syndrome : 0x08b3
                                | ({32{i_sel[640]}} & 32'h01000080)     //  syndrome : 0x12c9
                                | ({32{i_sel[639]}} & 32'h01000040)     //  syndrome : 0x0acc
                                | ({32{i_sel[638]}} & 32'h01000020)     //  syndrome : 0x06cf
                                | ({32{i_sel[637]}} & 32'h01000010)     //  syndrome : 0x15f7
                                | ({32{i_sel[636]}} & 32'h01000008)     //  syndrome : 0x1c6b
                                | ({32{i_sel[635]}} & 32'h01000004)     //  syndrome : 0x18a5
                                | ({32{i_sel[634]}} & 32'h01000002)     //  syndrome : 0x0ffa
                                | ({32{i_sel[633]}} & 32'h01000001)     //  syndrome : 0x116c
                                | ({32{i_sel[632]}} & 32'h01000000)     //  syndrome : 0x0b1f
                                | ({32{i_sel[631]}} & 32'h01000000)     //  syndrome : 0x131f
                                | ({32{i_sel[630]}} & 32'h01000000)     //  syndrome : 0x1f1f
                                | ({32{i_sel[629]}} & 32'h01000000)     //  syndrome : 0x191f
                                | ({32{i_sel[628]}} & 32'h01000000)     //  syndrome : 0x1a1f
                                | ({32{i_sel[627]}} & 32'h01000000)     //  syndrome : 0x1b9f
                                | ({32{i_sel[626]}} & 32'h01000000)     //  syndrome : 0x1b5f
                                | ({32{i_sel[625]}} & 32'h01000000)     //  syndrome : 0x1b3f
                                | ({32{i_sel[624]}} & 32'h01000000)     //  syndrome : 0x1b0f
                                | ({32{i_sel[623]}} & 32'h01000000)     //  syndrome : 0x1b17
                                | ({32{i_sel[622]}} & 32'h01000000)     //  syndrome : 0x1b1b
                                | ({32{i_sel[621]}} & 32'h01000000)     //  syndrome : 0x1b1d
                                | ({32{i_sel[620]}} & 32'h01000000)     //  syndrome : 0x1b1e
                                | ({32{i_sel[619]}} & 32'h00c00000)     //  syndrome : 0x01d5
                                | ({32{i_sel[618]}} & 32'h00a00000)     //  syndrome : 0x013e
                                | ({32{i_sel[617]}} & 32'h00900000)     //  syndrome : 0x1472
                                | ({32{i_sel[616]}} & 32'h00880000)     //  syndrome : 0x1ed4
                                | ({32{i_sel[615]}} & 32'h00840000)     //  syndrome : 0x0ebf
                                | ({32{i_sel[614]}} & 32'h00820000)     //  syndrome : 0x13b3
                                | ({32{i_sel[613]}} & 32'h00810000)     //  syndrome : 0x1d35
                                | ({32{i_sel[612]}} & 32'h00808000)     //  syndrome : 0x0f4e
                                | ({32{i_sel[611]}} & 32'h00804000)     //  syndrome : 0x134a
                                | ({32{i_sel[610]}} & 32'h00802000)     //  syndrome : 0x1d48
                                | ({32{i_sel[609]}} & 32'h00801000)     //  syndrome : 0x0f71
                                | ({32{i_sel[608]}} & 32'h00800800)     //  syndrome : 0x066c
                                | ({32{i_sel[607]}} & 32'h00800400)     //  syndrome : 0x02e3
                                | ({32{i_sel[606]}} & 32'h00800200)     //  syndrome : 0x159d
                                | ({32{i_sel[605]}} & 32'h00800100)     //  syndrome : 0x0b1a
                                | ({32{i_sel[604]}} & 32'h00800080)     //  syndrome : 0x1160
                                | ({32{i_sel[603]}} & 32'h00800040)     //  syndrome : 0x0965
                                | ({32{i_sel[602]}} & 32'h00800020)     //  syndrome : 0x0566
                                | ({32{i_sel[601]}} & 32'h00800010)     //  syndrome : 0x165e
                                | ({32{i_sel[600]}} & 32'h00800008)     //  syndrome : 0x1fc2
                                | ({32{i_sel[599]}} & 32'h00800004)     //  syndrome : 0x1b0c
                                | ({32{i_sel[598]}} & 32'h00800002)     //  syndrome : 0x0c53
                                | ({32{i_sel[597]}} & 32'h00800001)     //  syndrome : 0x12c5
                                | ({32{i_sel[596]}} & 32'h00800000)     //  syndrome : 0x08b6
                                | ({32{i_sel[595]}} & 32'h00800000)     //  syndrome : 0x10b6
                                | ({32{i_sel[594]}} & 32'h00800000)     //  syndrome : 0x1cb6
                                | ({32{i_sel[593]}} & 32'h00800000)     //  syndrome : 0x1ab6
                                | ({32{i_sel[592]}} & 32'h00800000)     //  syndrome : 0x19b6
                                | ({32{i_sel[591]}} & 32'h00800000)     //  syndrome : 0x1836
                                | ({32{i_sel[590]}} & 32'h00800000)     //  syndrome : 0x18f6
                                | ({32{i_sel[589]}} & 32'h00800000)     //  syndrome : 0x1896
                                | ({32{i_sel[588]}} & 32'h00800000)     //  syndrome : 0x18a6
                                | ({32{i_sel[587]}} & 32'h00800000)     //  syndrome : 0x18be
                                | ({32{i_sel[586]}} & 32'h00800000)     //  syndrome : 0x18b2
                                | ({32{i_sel[585]}} & 32'h00800000)     //  syndrome : 0x18b4
                                | ({32{i_sel[584]}} & 32'h00800000)     //  syndrome : 0x18b7
                                | ({32{i_sel[583]}} & 32'h00600000)     //  syndrome : 0x00eb
                                | ({32{i_sel[582]}} & 32'h00500000)     //  syndrome : 0x15a7
                                | ({32{i_sel[581]}} & 32'h00480000)     //  syndrome : 0x1f01
                                | ({32{i_sel[580]}} & 32'h00440000)     //  syndrome : 0x0f6a
                                | ({32{i_sel[579]}} & 32'h00420000)     //  syndrome : 0x1266
                                | ({32{i_sel[578]}} & 32'h00410000)     //  syndrome : 0x1ce0
                                | ({32{i_sel[577]}} & 32'h00408000)     //  syndrome : 0x0e9b
                                | ({32{i_sel[576]}} & 32'h00404000)     //  syndrome : 0x129f
                                | ({32{i_sel[575]}} & 32'h00402000)     //  syndrome : 0x1c9d
                                | ({32{i_sel[574]}} & 32'h00401000)     //  syndrome : 0x0ea4
                                | ({32{i_sel[573]}} & 32'h00400800)     //  syndrome : 0x07b9
                                | ({32{i_sel[572]}} & 32'h00400400)     //  syndrome : 0x0336
                                | ({32{i_sel[571]}} & 32'h00400200)     //  syndrome : 0x1448
                                | ({32{i_sel[570]}} & 32'h00400100)     //  syndrome : 0x0acf
                                | ({32{i_sel[569]}} & 32'h00400080)     //  syndrome : 0x10b5
                                | ({32{i_sel[568]}} & 32'h00400040)     //  syndrome : 0x08b0
                                | ({32{i_sel[567]}} & 32'h00400020)     //  syndrome : 0x04b3
                                | ({32{i_sel[566]}} & 32'h00400010)     //  syndrome : 0x178b
                                | ({32{i_sel[565]}} & 32'h00400008)     //  syndrome : 0x1e17
                                | ({32{i_sel[564]}} & 32'h00400004)     //  syndrome : 0x1ad9
                                | ({32{i_sel[563]}} & 32'h00400002)     //  syndrome : 0x0d86
                                | ({32{i_sel[562]}} & 32'h00400001)     //  syndrome : 0x1310
                                | ({32{i_sel[561]}} & 32'h00400000)     //  syndrome : 0x0963
                                | ({32{i_sel[560]}} & 32'h00400000)     //  syndrome : 0x1163
                                | ({32{i_sel[559]}} & 32'h00400000)     //  syndrome : 0x1d63
                                | ({32{i_sel[558]}} & 32'h00400000)     //  syndrome : 0x1b63
                                | ({32{i_sel[557]}} & 32'h00400000)     //  syndrome : 0x1863
                                | ({32{i_sel[556]}} & 32'h00400000)     //  syndrome : 0x19e3
                                | ({32{i_sel[555]}} & 32'h00400000)     //  syndrome : 0x1923
                                | ({32{i_sel[554]}} & 32'h00400000)     //  syndrome : 0x1943
                                | ({32{i_sel[553]}} & 32'h00400000)     //  syndrome : 0x1973
                                | ({32{i_sel[552]}} & 32'h00400000)     //  syndrome : 0x196b
                                | ({32{i_sel[551]}} & 32'h00400000)     //  syndrome : 0x1967
                                | ({32{i_sel[550]}} & 32'h00400000)     //  syndrome : 0x1961
                                | ({32{i_sel[549]}} & 32'h00400000)     //  syndrome : 0x1962
                                | ({32{i_sel[548]}} & 32'h00300000)     //  syndrome : 0x154c
                                | ({32{i_sel[547]}} & 32'h00280000)     //  syndrome : 0x1fea
                                | ({32{i_sel[546]}} & 32'h00240000)     //  syndrome : 0x0f81
                                | ({32{i_sel[545]}} & 32'h00220000)     //  syndrome : 0x128d
                                | ({32{i_sel[544]}} & 32'h00210000)     //  syndrome : 0x1c0b
                                | ({32{i_sel[543]}} & 32'h00208000)     //  syndrome : 0x0e70
                                | ({32{i_sel[542]}} & 32'h00204000)     //  syndrome : 0x1274
                                | ({32{i_sel[541]}} & 32'h00202000)     //  syndrome : 0x1c76
                                | ({32{i_sel[540]}} & 32'h00201000)     //  syndrome : 0x0e4f
                                | ({32{i_sel[539]}} & 32'h00200800)     //  syndrome : 0x0752
                                | ({32{i_sel[538]}} & 32'h00200400)     //  syndrome : 0x03dd
                                | ({32{i_sel[537]}} & 32'h00200200)     //  syndrome : 0x14a3
                                | ({32{i_sel[536]}} & 32'h00200100)     //  syndrome : 0x0a24
                                | ({32{i_sel[535]}} & 32'h00200080)     //  syndrome : 0x105e
                                | ({32{i_sel[534]}} & 32'h00200040)     //  syndrome : 0x085b
                                | ({32{i_sel[533]}} & 32'h00200020)     //  syndrome : 0x0458
                                | ({32{i_sel[532]}} & 32'h00200010)     //  syndrome : 0x1760
                                | ({32{i_sel[531]}} & 32'h00200008)     //  syndrome : 0x1efc
                                | ({32{i_sel[530]}} & 32'h00200004)     //  syndrome : 0x1a32
                                | ({32{i_sel[529]}} & 32'h00200002)     //  syndrome : 0x0d6d
                                | ({32{i_sel[528]}} & 32'h00200001)     //  syndrome : 0x13fb
                                | ({32{i_sel[527]}} & 32'h00200000)     //  syndrome : 0x0988
                                | ({32{i_sel[526]}} & 32'h00200000)     //  syndrome : 0x1188
                                | ({32{i_sel[525]}} & 32'h00200000)     //  syndrome : 0x1d88
                                | ({32{i_sel[524]}} & 32'h00200000)     //  syndrome : 0x1b88
                                | ({32{i_sel[523]}} & 32'h00200000)     //  syndrome : 0x1888
                                | ({32{i_sel[522]}} & 32'h00200000)     //  syndrome : 0x1908
                                | ({32{i_sel[521]}} & 32'h00200000)     //  syndrome : 0x19c8
                                | ({32{i_sel[520]}} & 32'h00200000)     //  syndrome : 0x19a8
                                | ({32{i_sel[519]}} & 32'h00200000)     //  syndrome : 0x1998
                                | ({32{i_sel[518]}} & 32'h00200000)     //  syndrome : 0x1980
                                | ({32{i_sel[517]}} & 32'h00200000)     //  syndrome : 0x198c
                                | ({32{i_sel[516]}} & 32'h00200000)     //  syndrome : 0x198a
                                | ({32{i_sel[515]}} & 32'h00200000)     //  syndrome : 0x1989
                                | ({32{i_sel[514]}} & 32'h00180000)     //  syndrome : 0x0aa6
                                | ({32{i_sel[513]}} & 32'h00140000)     //  syndrome : 0x1acd
                                | ({32{i_sel[512]}} & 32'h00120000)     //  syndrome : 0x07c1
                                | ({32{i_sel[511]}} & 32'h00110000)     //  syndrome : 0x0947
                                | ({32{i_sel[510]}} & 32'h00108000)     //  syndrome : 0x1b3c
                                | ({32{i_sel[509]}} & 32'h00104000)     //  syndrome : 0x0738
                                | ({32{i_sel[508]}} & 32'h00102000)     //  syndrome : 0x093a
                                | ({32{i_sel[507]}} & 32'h00101000)     //  syndrome : 0x1b03
                                | ({32{i_sel[506]}} & 32'h00100800)     //  syndrome : 0x121e
                                | ({32{i_sel[505]}} & 32'h00100400)     //  syndrome : 0x1691
                                | ({32{i_sel[504]}} & 32'h00100200)     //  syndrome : 0x01ef
                                | ({32{i_sel[503]}} & 32'h00100100)     //  syndrome : 0x1f68
                                | ({32{i_sel[502]}} & 32'h00100080)     //  syndrome : 0x0512
                                | ({32{i_sel[501]}} & 32'h00100040)     //  syndrome : 0x1d17
                                | ({32{i_sel[500]}} & 32'h00100020)     //  syndrome : 0x1114
                                | ({32{i_sel[499]}} & 32'h00100010)     //  syndrome : 0x022c
                                | ({32{i_sel[498]}} & 32'h00100008)     //  syndrome : 0x0bb0
                                | ({32{i_sel[497]}} & 32'h00100004)     //  syndrome : 0x0f7e
                                | ({32{i_sel[496]}} & 32'h00100002)     //  syndrome : 0x1821
                                | ({32{i_sel[495]}} & 32'h00100001)     //  syndrome : 0x06b7
                                | ({32{i_sel[494]}} & 32'h00100000)     //  syndrome : 0x1cc4
                                | ({32{i_sel[493]}} & 32'h00100000)     //  syndrome : 0x04c4
                                | ({32{i_sel[492]}} & 32'h00100000)     //  syndrome : 0x08c4
                                | ({32{i_sel[491]}} & 32'h00100000)     //  syndrome : 0x0ec4
                                | ({32{i_sel[490]}} & 32'h00100000)     //  syndrome : 0x0dc4
                                | ({32{i_sel[489]}} & 32'h00100000)     //  syndrome : 0x0c44
                                | ({32{i_sel[488]}} & 32'h00100000)     //  syndrome : 0x0c84
                                | ({32{i_sel[487]}} & 32'h00100000)     //  syndrome : 0x0ce4
                                | ({32{i_sel[486]}} & 32'h00100000)     //  syndrome : 0x0cd4
                                | ({32{i_sel[485]}} & 32'h00100000)     //  syndrome : 0x0ccc
                                | ({32{i_sel[484]}} & 32'h00100000)     //  syndrome : 0x0cc0
                                | ({32{i_sel[483]}} & 32'h00100000)     //  syndrome : 0x0cc6
                                | ({32{i_sel[482]}} & 32'h00100000)     //  syndrome : 0x0cc5
                                | ({32{i_sel[481]}} & 32'h000c0000)     //  syndrome : 0x106b
                                | ({32{i_sel[480]}} & 32'h000a0000)     //  syndrome : 0x0d67
                                | ({32{i_sel[479]}} & 32'h00090000)     //  syndrome : 0x03e1
                                | ({32{i_sel[478]}} & 32'h00088000)     //  syndrome : 0x119a
                                | ({32{i_sel[477]}} & 32'h00084000)     //  syndrome : 0x0d9e
                                | ({32{i_sel[476]}} & 32'h00082000)     //  syndrome : 0x039c
                                | ({32{i_sel[475]}} & 32'h00081000)     //  syndrome : 0x11a5
                                | ({32{i_sel[474]}} & 32'h00080800)     //  syndrome : 0x18b8
                                | ({32{i_sel[473]}} & 32'h00080400)     //  syndrome : 0x1c37
                                | ({32{i_sel[472]}} & 32'h00080200)     //  syndrome : 0x0b49
                                | ({32{i_sel[471]}} & 32'h00080100)     //  syndrome : 0x15ce
                                | ({32{i_sel[470]}} & 32'h00080080)     //  syndrome : 0x0fb4
                                | ({32{i_sel[469]}} & 32'h00080040)     //  syndrome : 0x17b1
                                | ({32{i_sel[468]}} & 32'h00080020)     //  syndrome : 0x1bb2
                                | ({32{i_sel[467]}} & 32'h00080010)     //  syndrome : 0x088a
                                | ({32{i_sel[466]}} & 32'h00080008)     //  syndrome : 0x0116
                                | ({32{i_sel[465]}} & 32'h00080004)     //  syndrome : 0x05d8
                                | ({32{i_sel[464]}} & 32'h00080002)     //  syndrome : 0x1287
                                | ({32{i_sel[463]}} & 32'h00080001)     //  syndrome : 0x0c11
                                | ({32{i_sel[462]}} & 32'h00080000)     //  syndrome : 0x1662
                                | ({32{i_sel[461]}} & 32'h00080000)     //  syndrome : 0x0e62
                                | ({32{i_sel[460]}} & 32'h00080000)     //  syndrome : 0x0262
                                | ({32{i_sel[459]}} & 32'h00080000)     //  syndrome : 0x0462
                                | ({32{i_sel[458]}} & 32'h00080000)     //  syndrome : 0x0762
                                | ({32{i_sel[457]}} & 32'h00080000)     //  syndrome : 0x06e2
                                | ({32{i_sel[456]}} & 32'h00080000)     //  syndrome : 0x0622
                                | ({32{i_sel[455]}} & 32'h00080000)     //  syndrome : 0x0642
                                | ({32{i_sel[454]}} & 32'h00080000)     //  syndrome : 0x0672
                                | ({32{i_sel[453]}} & 32'h00080000)     //  syndrome : 0x066a
                                | ({32{i_sel[452]}} & 32'h00080000)     //  syndrome : 0x0666
                                | ({32{i_sel[451]}} & 32'h00080000)     //  syndrome : 0x0660
                                | ({32{i_sel[450]}} & 32'h00080000)     //  syndrome : 0x0663
                                | ({32{i_sel[449]}} & 32'h00060000)     //  syndrome : 0x1d0c
                                | ({32{i_sel[448]}} & 32'h00050000)     //  syndrome : 0x138a
                                | ({32{i_sel[447]}} & 32'h00048000)     //  syndrome : 0x01f1
                                | ({32{i_sel[446]}} & 32'h00044000)     //  syndrome : 0x1df5
                                | ({32{i_sel[445]}} & 32'h00042000)     //  syndrome : 0x13f7
                                | ({32{i_sel[444]}} & 32'h00041000)     //  syndrome : 0x01ce
                                | ({32{i_sel[443]}} & 32'h00040800)     //  syndrome : 0x08d3
                                | ({32{i_sel[442]}} & 32'h00040400)     //  syndrome : 0x0c5c
                                | ({32{i_sel[441]}} & 32'h00040200)     //  syndrome : 0x1b22
                                | ({32{i_sel[440]}} & 32'h00040100)     //  syndrome : 0x05a5
                                | ({32{i_sel[439]}} & 32'h00040080)     //  syndrome : 0x1fdf
                                | ({32{i_sel[438]}} & 32'h00040040)     //  syndrome : 0x07da
                                | ({32{i_sel[437]}} & 32'h00040020)     //  syndrome : 0x0bd9
                                | ({32{i_sel[436]}} & 32'h00040010)     //  syndrome : 0x18e1
                                | ({32{i_sel[435]}} & 32'h00040008)     //  syndrome : 0x117d
                                | ({32{i_sel[434]}} & 32'h00040004)     //  syndrome : 0x15b3
                                | ({32{i_sel[433]}} & 32'h00040002)     //  syndrome : 0x02ec
                                | ({32{i_sel[432]}} & 32'h00040001)     //  syndrome : 0x1c7a
                                | ({32{i_sel[431]}} & 32'h00040000)     //  syndrome : 0x0609
                                | ({32{i_sel[430]}} & 32'h00040000)     //  syndrome : 0x1e09
                                | ({32{i_sel[429]}} & 32'h00040000)     //  syndrome : 0x1209
                                | ({32{i_sel[428]}} & 32'h00040000)     //  syndrome : 0x1409
                                | ({32{i_sel[427]}} & 32'h00040000)     //  syndrome : 0x1709
                                | ({32{i_sel[426]}} & 32'h00040000)     //  syndrome : 0x1689
                                | ({32{i_sel[425]}} & 32'h00040000)     //  syndrome : 0x1649
                                | ({32{i_sel[424]}} & 32'h00040000)     //  syndrome : 0x1629
                                | ({32{i_sel[423]}} & 32'h00040000)     //  syndrome : 0x1619
                                | ({32{i_sel[422]}} & 32'h00040000)     //  syndrome : 0x1601
                                | ({32{i_sel[421]}} & 32'h00040000)     //  syndrome : 0x160d
                                | ({32{i_sel[420]}} & 32'h00040000)     //  syndrome : 0x160b
                                | ({32{i_sel[419]}} & 32'h00040000)     //  syndrome : 0x1608
                                | ({32{i_sel[418]}} & 32'h00030000)     //  syndrome : 0x0e86
                                | ({32{i_sel[417]}} & 32'h00028000)     //  syndrome : 0x1cfd
                                | ({32{i_sel[416]}} & 32'h00024000)     //  syndrome : 0x00f9
                                | ({32{i_sel[415]}} & 32'h00022000)     //  syndrome : 0x0efb
                                | ({32{i_sel[414]}} & 32'h00021000)     //  syndrome : 0x1cc2
                                | ({32{i_sel[413]}} & 32'h00020800)     //  syndrome : 0x15df
                                | ({32{i_sel[412]}} & 32'h00020400)     //  syndrome : 0x1150
                                | ({32{i_sel[411]}} & 32'h00020200)     //  syndrome : 0x062e
                                | ({32{i_sel[410]}} & 32'h00020100)     //  syndrome : 0x18a9
                                | ({32{i_sel[409]}} & 32'h00020080)     //  syndrome : 0x02d3
                                | ({32{i_sel[408]}} & 32'h00020040)     //  syndrome : 0x1ad6
                                | ({32{i_sel[407]}} & 32'h00020020)     //  syndrome : 0x16d5
                                | ({32{i_sel[406]}} & 32'h00020010)     //  syndrome : 0x05ed
                                | ({32{i_sel[405]}} & 32'h00020008)     //  syndrome : 0x0c71
                                | ({32{i_sel[404]}} & 32'h00020004)     //  syndrome : 0x08bf
                                | ({32{i_sel[403]}} & 32'h00020002)     //  syndrome : 0x1fe0
                                | ({32{i_sel[402]}} & 32'h00020001)     //  syndrome : 0x0176
                                | ({32{i_sel[401]}} & 32'h00020000)     //  syndrome : 0x1b05
                                | ({32{i_sel[400]}} & 32'h00020000)     //  syndrome : 0x0305
                                | ({32{i_sel[399]}} & 32'h00020000)     //  syndrome : 0x0f05
                                | ({32{i_sel[398]}} & 32'h00020000)     //  syndrome : 0x0905
                                | ({32{i_sel[397]}} & 32'h00020000)     //  syndrome : 0x0a05
                                | ({32{i_sel[396]}} & 32'h00020000)     //  syndrome : 0x0b85
                                | ({32{i_sel[395]}} & 32'h00020000)     //  syndrome : 0x0b45
                                | ({32{i_sel[394]}} & 32'h00020000)     //  syndrome : 0x0b25
                                | ({32{i_sel[393]}} & 32'h00020000)     //  syndrome : 0x0b15
                                | ({32{i_sel[392]}} & 32'h00020000)     //  syndrome : 0x0b0d
                                | ({32{i_sel[391]}} & 32'h00020000)     //  syndrome : 0x0b01
                                | ({32{i_sel[390]}} & 32'h00020000)     //  syndrome : 0x0b07
                                | ({32{i_sel[389]}} & 32'h00020000)     //  syndrome : 0x0b04
                                | ({32{i_sel[388]}} & 32'h00018000)     //  syndrome : 0x127b
                                | ({32{i_sel[387]}} & 32'h00014000)     //  syndrome : 0x0e7f
                                | ({32{i_sel[386]}} & 32'h00012000)     //  syndrome : 0x007d
                                | ({32{i_sel[385]}} & 32'h00011000)     //  syndrome : 0x1244
                                | ({32{i_sel[384]}} & 32'h00010800)     //  syndrome : 0x1b59
                                | ({32{i_sel[383]}} & 32'h00010400)     //  syndrome : 0x1fd6
                                | ({32{i_sel[382]}} & 32'h00010200)     //  syndrome : 0x08a8
                                | ({32{i_sel[381]}} & 32'h00010100)     //  syndrome : 0x162f
                                | ({32{i_sel[380]}} & 32'h00010080)     //  syndrome : 0x0c55
                                | ({32{i_sel[379]}} & 32'h00010040)     //  syndrome : 0x1450
                                | ({32{i_sel[378]}} & 32'h00010020)     //  syndrome : 0x1853
                                | ({32{i_sel[377]}} & 32'h00010010)     //  syndrome : 0x0b6b
                                | ({32{i_sel[376]}} & 32'h00010008)     //  syndrome : 0x02f7
                                | ({32{i_sel[375]}} & 32'h00010004)     //  syndrome : 0x0639
                                | ({32{i_sel[374]}} & 32'h00010002)     //  syndrome : 0x1166
                                | ({32{i_sel[373]}} & 32'h00010001)     //  syndrome : 0x0ff0
                                | ({32{i_sel[372]}} & 32'h00010000)     //  syndrome : 0x1583
                                | ({32{i_sel[371]}} & 32'h00010000)     //  syndrome : 0x0d83
                                | ({32{i_sel[370]}} & 32'h00010000)     //  syndrome : 0x0183
                                | ({32{i_sel[369]}} & 32'h00010000)     //  syndrome : 0x0783
                                | ({32{i_sel[368]}} & 32'h00010000)     //  syndrome : 0x0483
                                | ({32{i_sel[367]}} & 32'h00010000)     //  syndrome : 0x0503
                                | ({32{i_sel[366]}} & 32'h00010000)     //  syndrome : 0x05c3
                                | ({32{i_sel[365]}} & 32'h00010000)     //  syndrome : 0x05a3
                                | ({32{i_sel[364]}} & 32'h00010000)     //  syndrome : 0x0593
                                | ({32{i_sel[363]}} & 32'h00010000)     //  syndrome : 0x058b
                                | ({32{i_sel[362]}} & 32'h00010000)     //  syndrome : 0x0587
                                | ({32{i_sel[361]}} & 32'h00010000)     //  syndrome : 0x0581
                                | ({32{i_sel[360]}} & 32'h00010000)     //  syndrome : 0x0582
                                | ({32{i_sel[359]}} & 32'h0000c000)     //  syndrome : 0x1c04
                                | ({32{i_sel[358]}} & 32'h0000a000)     //  syndrome : 0x1206
                                | ({32{i_sel[357]}} & 32'h00009000)     //  syndrome : 0x003f
                                | ({32{i_sel[356]}} & 32'h00008800)     //  syndrome : 0x0922
                                | ({32{i_sel[355]}} & 32'h00008400)     //  syndrome : 0x0dad
                                | ({32{i_sel[354]}} & 32'h00008200)     //  syndrome : 0x1ad3
                                | ({32{i_sel[353]}} & 32'h00008100)     //  syndrome : 0x0454
                                | ({32{i_sel[352]}} & 32'h00008080)     //  syndrome : 0x1e2e
                                | ({32{i_sel[351]}} & 32'h00008040)     //  syndrome : 0x062b
                                | ({32{i_sel[350]}} & 32'h00008020)     //  syndrome : 0x0a28
                                | ({32{i_sel[349]}} & 32'h00008010)     //  syndrome : 0x1910
                                | ({32{i_sel[348]}} & 32'h00008008)     //  syndrome : 0x108c
                                | ({32{i_sel[347]}} & 32'h00008004)     //  syndrome : 0x1442
                                | ({32{i_sel[346]}} & 32'h00008002)     //  syndrome : 0x031d
                                | ({32{i_sel[345]}} & 32'h00008001)     //  syndrome : 0x1d8b
                                | ({32{i_sel[344]}} & 32'h00008000)     //  syndrome : 0x07f8
                                | ({32{i_sel[343]}} & 32'h00008000)     //  syndrome : 0x1ff8
                                | ({32{i_sel[342]}} & 32'h00008000)     //  syndrome : 0x13f8
                                | ({32{i_sel[341]}} & 32'h00008000)     //  syndrome : 0x15f8
                                | ({32{i_sel[340]}} & 32'h00008000)     //  syndrome : 0x16f8
                                | ({32{i_sel[339]}} & 32'h00008000)     //  syndrome : 0x1778
                                | ({32{i_sel[338]}} & 32'h00008000)     //  syndrome : 0x17b8
                                | ({32{i_sel[337]}} & 32'h00008000)     //  syndrome : 0x17d8
                                | ({32{i_sel[336]}} & 32'h00008000)     //  syndrome : 0x17e8
                                | ({32{i_sel[335]}} & 32'h00008000)     //  syndrome : 0x17f0
                                | ({32{i_sel[334]}} & 32'h00008000)     //  syndrome : 0x17fc
                                | ({32{i_sel[333]}} & 32'h00008000)     //  syndrome : 0x17fa
                                | ({32{i_sel[332]}} & 32'h00008000)     //  syndrome : 0x17f9
                                | ({32{i_sel[331]}} & 32'h00006000)     //  syndrome : 0x0e02
                                | ({32{i_sel[330]}} & 32'h00005000)     //  syndrome : 0x1c3b
                                | ({32{i_sel[329]}} & 32'h00004800)     //  syndrome : 0x1526
                                | ({32{i_sel[328]}} & 32'h00004400)     //  syndrome : 0x11a9
                                | ({32{i_sel[327]}} & 32'h00004200)     //  syndrome : 0x06d7
                                | ({32{i_sel[326]}} & 32'h00004100)     //  syndrome : 0x1850
                                | ({32{i_sel[325]}} & 32'h00004080)     //  syndrome : 0x022a
                                | ({32{i_sel[324]}} & 32'h00004040)     //  syndrome : 0x1a2f
                                | ({32{i_sel[323]}} & 32'h00004020)     //  syndrome : 0x162c
                                | ({32{i_sel[322]}} & 32'h00004010)     //  syndrome : 0x0514
                                | ({32{i_sel[321]}} & 32'h00004008)     //  syndrome : 0x0c88
                                | ({32{i_sel[320]}} & 32'h00004004)     //  syndrome : 0x0846
                                | ({32{i_sel[319]}} & 32'h00004002)     //  syndrome : 0x1f19
                                | ({32{i_sel[318]}} & 32'h00004001)     //  syndrome : 0x018f
                                | ({32{i_sel[317]}} & 32'h00004000)     //  syndrome : 0x1bfc
                                | ({32{i_sel[316]}} & 32'h00004000)     //  syndrome : 0x03fc
                                | ({32{i_sel[315]}} & 32'h00004000)     //  syndrome : 0x0ffc
                                | ({32{i_sel[314]}} & 32'h00004000)     //  syndrome : 0x09fc
                                | ({32{i_sel[313]}} & 32'h00004000)     //  syndrome : 0x0afc
                                | ({32{i_sel[312]}} & 32'h00004000)     //  syndrome : 0x0b7c
                                | ({32{i_sel[311]}} & 32'h00004000)     //  syndrome : 0x0bbc
                                | ({32{i_sel[310]}} & 32'h00004000)     //  syndrome : 0x0bdc
                                | ({32{i_sel[309]}} & 32'h00004000)     //  syndrome : 0x0bec
                                | ({32{i_sel[308]}} & 32'h00004000)     //  syndrome : 0x0bf4
                                | ({32{i_sel[307]}} & 32'h00004000)     //  syndrome : 0x0bf8
                                | ({32{i_sel[306]}} & 32'h00004000)     //  syndrome : 0x0bfe
                                | ({32{i_sel[305]}} & 32'h00004000)     //  syndrome : 0x0bfd
                                | ({32{i_sel[304]}} & 32'h00003000)     //  syndrome : 0x1239
                                | ({32{i_sel[303]}} & 32'h00002800)     //  syndrome : 0x1b24
                                | ({32{i_sel[302]}} & 32'h00002400)     //  syndrome : 0x1fab
                                | ({32{i_sel[301]}} & 32'h00002200)     //  syndrome : 0x08d5
                                | ({32{i_sel[300]}} & 32'h00002100)     //  syndrome : 0x1652
                                | ({32{i_sel[299]}} & 32'h00002080)     //  syndrome : 0x0c28
                                | ({32{i_sel[298]}} & 32'h00002040)     //  syndrome : 0x142d
                                | ({32{i_sel[297]}} & 32'h00002020)     //  syndrome : 0x182e
                                | ({32{i_sel[296]}} & 32'h00002010)     //  syndrome : 0x0b16
                                | ({32{i_sel[295]}} & 32'h00002008)     //  syndrome : 0x028a
                                | ({32{i_sel[294]}} & 32'h00002004)     //  syndrome : 0x0644
                                | ({32{i_sel[293]}} & 32'h00002002)     //  syndrome : 0x111b
                                | ({32{i_sel[292]}} & 32'h00002001)     //  syndrome : 0x0f8d
                                | ({32{i_sel[291]}} & 32'h00002000)     //  syndrome : 0x15fe
                                | ({32{i_sel[290]}} & 32'h00002000)     //  syndrome : 0x0dfe
                                | ({32{i_sel[289]}} & 32'h00002000)     //  syndrome : 0x01fe
                                | ({32{i_sel[288]}} & 32'h00002000)     //  syndrome : 0x07fe
                                | ({32{i_sel[287]}} & 32'h00002000)     //  syndrome : 0x04fe
                                | ({32{i_sel[286]}} & 32'h00002000)     //  syndrome : 0x057e
                                | ({32{i_sel[285]}} & 32'h00002000)     //  syndrome : 0x05be
                                | ({32{i_sel[284]}} & 32'h00002000)     //  syndrome : 0x05de
                                | ({32{i_sel[283]}} & 32'h00002000)     //  syndrome : 0x05ee
                                | ({32{i_sel[282]}} & 32'h00002000)     //  syndrome : 0x05f6
                                | ({32{i_sel[281]}} & 32'h00002000)     //  syndrome : 0x05fa
                                | ({32{i_sel[280]}} & 32'h00002000)     //  syndrome : 0x05fc
                                | ({32{i_sel[279]}} & 32'h00002000)     //  syndrome : 0x05ff
                                | ({32{i_sel[278]}} & 32'h00001800)     //  syndrome : 0x091d
                                | ({32{i_sel[277]}} & 32'h00001400)     //  syndrome : 0x0d92
                                | ({32{i_sel[276]}} & 32'h00001200)     //  syndrome : 0x1aec
                                | ({32{i_sel[275]}} & 32'h00001100)     //  syndrome : 0x046b
                                | ({32{i_sel[274]}} & 32'h00001080)     //  syndrome : 0x1e11
                                | ({32{i_sel[273]}} & 32'h00001040)     //  syndrome : 0x0614
                                | ({32{i_sel[272]}} & 32'h00001020)     //  syndrome : 0x0a17
                                | ({32{i_sel[271]}} & 32'h00001010)     //  syndrome : 0x192f
                                | ({32{i_sel[270]}} & 32'h00001008)     //  syndrome : 0x10b3
                                | ({32{i_sel[269]}} & 32'h00001004)     //  syndrome : 0x147d
                                | ({32{i_sel[268]}} & 32'h00001002)     //  syndrome : 0x0322
                                | ({32{i_sel[267]}} & 32'h00001001)     //  syndrome : 0x1db4
                                | ({32{i_sel[266]}} & 32'h00001000)     //  syndrome : 0x07c7
                                | ({32{i_sel[265]}} & 32'h00001000)     //  syndrome : 0x1fc7
                                | ({32{i_sel[264]}} & 32'h00001000)     //  syndrome : 0x13c7
                                | ({32{i_sel[263]}} & 32'h00001000)     //  syndrome : 0x15c7
                                | ({32{i_sel[262]}} & 32'h00001000)     //  syndrome : 0x16c7
                                | ({32{i_sel[261]}} & 32'h00001000)     //  syndrome : 0x1747
                                | ({32{i_sel[260]}} & 32'h00001000)     //  syndrome : 0x1787
                                | ({32{i_sel[259]}} & 32'h00001000)     //  syndrome : 0x17e7
                                | ({32{i_sel[258]}} & 32'h00001000)     //  syndrome : 0x17d7
                                | ({32{i_sel[257]}} & 32'h00001000)     //  syndrome : 0x17cf
                                | ({32{i_sel[256]}} & 32'h00001000)     //  syndrome : 0x17c3
                                | ({32{i_sel[255]}} & 32'h00001000)     //  syndrome : 0x17c5
                                | ({32{i_sel[254]}} & 32'h00001000)     //  syndrome : 0x17c6
                                | ({32{i_sel[253]}} & 32'h00000c00)     //  syndrome : 0x048f
                                | ({32{i_sel[252]}} & 32'h00000a00)     //  syndrome : 0x13f1
                                | ({32{i_sel[251]}} & 32'h00000900)     //  syndrome : 0x0d76
                                | ({32{i_sel[250]}} & 32'h00000880)     //  syndrome : 0x170c
                                | ({32{i_sel[249]}} & 32'h00000840)     //  syndrome : 0x0f09
                                | ({32{i_sel[248]}} & 32'h00000820)     //  syndrome : 0x030a
                                | ({32{i_sel[247]}} & 32'h00000810)     //  syndrome : 0x1032
                                | ({32{i_sel[246]}} & 32'h00000808)     //  syndrome : 0x19ae
                                | ({32{i_sel[245]}} & 32'h00000804)     //  syndrome : 0x1d60
                                | ({32{i_sel[244]}} & 32'h00000802)     //  syndrome : 0x0a3f
                                | ({32{i_sel[243]}} & 32'h00000801)     //  syndrome : 0x14a9
                                | ({32{i_sel[242]}} & 32'h00000800)     //  syndrome : 0x0eda
                                | ({32{i_sel[241]}} & 32'h00000800)     //  syndrome : 0x16da
                                | ({32{i_sel[240]}} & 32'h00000800)     //  syndrome : 0x1ada
                                | ({32{i_sel[239]}} & 32'h00000800)     //  syndrome : 0x1cda
                                | ({32{i_sel[238]}} & 32'h00000800)     //  syndrome : 0x1fda
                                | ({32{i_sel[237]}} & 32'h00000800)     //  syndrome : 0x1e5a
                                | ({32{i_sel[236]}} & 32'h00000800)     //  syndrome : 0x1e9a
                                | ({32{i_sel[235]}} & 32'h00000800)     //  syndrome : 0x1efa
                                | ({32{i_sel[234]}} & 32'h00000800)     //  syndrome : 0x1eca
                                | ({32{i_sel[233]}} & 32'h00000800)     //  syndrome : 0x1ed2
                                | ({32{i_sel[232]}} & 32'h00000800)     //  syndrome : 0x1ede
                                | ({32{i_sel[231]}} & 32'h00000800)     //  syndrome : 0x1ed8
                                | ({32{i_sel[230]}} & 32'h00000800)     //  syndrome : 0x1edb
                                | ({32{i_sel[229]}} & 32'h00000600)     //  syndrome : 0x177e
                                | ({32{i_sel[228]}} & 32'h00000500)     //  syndrome : 0x09f9
                                | ({32{i_sel[227]}} & 32'h00000480)     //  syndrome : 0x1383
                                | ({32{i_sel[226]}} & 32'h00000440)     //  syndrome : 0x0b86
                                | ({32{i_sel[225]}} & 32'h00000420)     //  syndrome : 0x0785
                                | ({32{i_sel[224]}} & 32'h00000410)     //  syndrome : 0x14bd
                                | ({32{i_sel[223]}} & 32'h00000408)     //  syndrome : 0x1d21
                                | ({32{i_sel[222]}} & 32'h00000404)     //  syndrome : 0x19ef
                                | ({32{i_sel[221]}} & 32'h00000402)     //  syndrome : 0x0eb0
                                | ({32{i_sel[220]}} & 32'h00000401)     //  syndrome : 0x1026
                                | ({32{i_sel[219]}} & 32'h00000400)     //  syndrome : 0x0a55
                                | ({32{i_sel[218]}} & 32'h00000400)     //  syndrome : 0x1255
                                | ({32{i_sel[217]}} & 32'h00000400)     //  syndrome : 0x1e55
                                | ({32{i_sel[216]}} & 32'h00000400)     //  syndrome : 0x1855
                                | ({32{i_sel[215]}} & 32'h00000400)     //  syndrome : 0x1b55
                                | ({32{i_sel[214]}} & 32'h00000400)     //  syndrome : 0x1ad5
                                | ({32{i_sel[213]}} & 32'h00000400)     //  syndrome : 0x1a15
                                | ({32{i_sel[212]}} & 32'h00000400)     //  syndrome : 0x1a75
                                | ({32{i_sel[211]}} & 32'h00000400)     //  syndrome : 0x1a45
                                | ({32{i_sel[210]}} & 32'h00000400)     //  syndrome : 0x1a5d
                                | ({32{i_sel[209]}} & 32'h00000400)     //  syndrome : 0x1a51
                                | ({32{i_sel[208]}} & 32'h00000400)     //  syndrome : 0x1a57
                                | ({32{i_sel[207]}} & 32'h00000400)     //  syndrome : 0x1a54
                                | ({32{i_sel[206]}} & 32'h00000300)     //  syndrome : 0x1e87
                                | ({32{i_sel[205]}} & 32'h00000280)     //  syndrome : 0x04fd
                                | ({32{i_sel[204]}} & 32'h00000240)     //  syndrome : 0x1cf8
                                | ({32{i_sel[203]}} & 32'h00000220)     //  syndrome : 0x10fb
                                | ({32{i_sel[202]}} & 32'h00000210)     //  syndrome : 0x03c3
                                | ({32{i_sel[201]}} & 32'h00000208)     //  syndrome : 0x0a5f
                                | ({32{i_sel[200]}} & 32'h00000204)     //  syndrome : 0x0e91
                                | ({32{i_sel[199]}} & 32'h00000202)     //  syndrome : 0x19ce
                                | ({32{i_sel[198]}} & 32'h00000201)     //  syndrome : 0x0758
                                | ({32{i_sel[197]}} & 32'h00000200)     //  syndrome : 0x1d2b
                                | ({32{i_sel[196]}} & 32'h00000200)     //  syndrome : 0x052b
                                | ({32{i_sel[195]}} & 32'h00000200)     //  syndrome : 0x092b
                                | ({32{i_sel[194]}} & 32'h00000200)     //  syndrome : 0x0f2b
                                | ({32{i_sel[193]}} & 32'h00000200)     //  syndrome : 0x0c2b
                                | ({32{i_sel[192]}} & 32'h00000200)     //  syndrome : 0x0dab
                                | ({32{i_sel[191]}} & 32'h00000200)     //  syndrome : 0x0d6b
                                | ({32{i_sel[190]}} & 32'h00000200)     //  syndrome : 0x0d0b
                                | ({32{i_sel[189]}} & 32'h00000200)     //  syndrome : 0x0d3b
                                | ({32{i_sel[188]}} & 32'h00000200)     //  syndrome : 0x0d23
                                | ({32{i_sel[187]}} & 32'h00000200)     //  syndrome : 0x0d2f
                                | ({32{i_sel[186]}} & 32'h00000200)     //  syndrome : 0x0d29
                                | ({32{i_sel[185]}} & 32'h00000200)     //  syndrome : 0x0d2a
                                | ({32{i_sel[184]}} & 32'h00000180)     //  syndrome : 0x1a7a
                                | ({32{i_sel[183]}} & 32'h00000140)     //  syndrome : 0x027f
                                | ({32{i_sel[182]}} & 32'h00000120)     //  syndrome : 0x0e7c
                                | ({32{i_sel[181]}} & 32'h00000110)     //  syndrome : 0x1d44
                                | ({32{i_sel[180]}} & 32'h00000108)     //  syndrome : 0x14d8
                                | ({32{i_sel[179]}} & 32'h00000104)     //  syndrome : 0x1016
                                | ({32{i_sel[178]}} & 32'h00000102)     //  syndrome : 0x0749
                                | ({32{i_sel[177]}} & 32'h00000101)     //  syndrome : 0x19df
                                | ({32{i_sel[176]}} & 32'h00000100)     //  syndrome : 0x03ac
                                | ({32{i_sel[175]}} & 32'h00000100)     //  syndrome : 0x1bac
                                | ({32{i_sel[174]}} & 32'h00000100)     //  syndrome : 0x17ac
                                | ({32{i_sel[173]}} & 32'h00000100)     //  syndrome : 0x11ac
                                | ({32{i_sel[172]}} & 32'h00000100)     //  syndrome : 0x12ac
                                | ({32{i_sel[171]}} & 32'h00000100)     //  syndrome : 0x132c
                                | ({32{i_sel[170]}} & 32'h00000100)     //  syndrome : 0x13ec
                                | ({32{i_sel[169]}} & 32'h00000100)     //  syndrome : 0x138c
                                | ({32{i_sel[168]}} & 32'h00000100)     //  syndrome : 0x13bc
                                | ({32{i_sel[167]}} & 32'h00000100)     //  syndrome : 0x13a4
                                | ({32{i_sel[166]}} & 32'h00000100)     //  syndrome : 0x13a8
                                | ({32{i_sel[165]}} & 32'h00000100)     //  syndrome : 0x13ae
                                | ({32{i_sel[164]}} & 32'h00000100)     //  syndrome : 0x13ad
                                | ({32{i_sel[163]}} & 32'h000000c0)     //  syndrome : 0x1805
                                | ({32{i_sel[162]}} & 32'h000000a0)     //  syndrome : 0x1406
                                | ({32{i_sel[161]}} & 32'h00000090)     //  syndrome : 0x073e
                                | ({32{i_sel[160]}} & 32'h00000088)     //  syndrome : 0x0ea2
                                | ({32{i_sel[159]}} & 32'h00000084)     //  syndrome : 0x0a6c
                                | ({32{i_sel[158]}} & 32'h00000082)     //  syndrome : 0x1d33
                                | ({32{i_sel[157]}} & 32'h00000081)     //  syndrome : 0x03a5
                                | ({32{i_sel[156]}} & 32'h00000080)     //  syndrome : 0x19d6
                                | ({32{i_sel[155]}} & 32'h00000080)     //  syndrome : 0x01d6
                                | ({32{i_sel[154]}} & 32'h00000080)     //  syndrome : 0x0dd6
                                | ({32{i_sel[153]}} & 32'h00000080)     //  syndrome : 0x0bd6
                                | ({32{i_sel[152]}} & 32'h00000080)     //  syndrome : 0x08d6
                                | ({32{i_sel[151]}} & 32'h00000080)     //  syndrome : 0x0956
                                | ({32{i_sel[150]}} & 32'h00000080)     //  syndrome : 0x0996
                                | ({32{i_sel[149]}} & 32'h00000080)     //  syndrome : 0x09f6
                                | ({32{i_sel[148]}} & 32'h00000080)     //  syndrome : 0x09c6
                                | ({32{i_sel[147]}} & 32'h00000080)     //  syndrome : 0x09de
                                | ({32{i_sel[146]}} & 32'h00000080)     //  syndrome : 0x09d2
                                | ({32{i_sel[145]}} & 32'h00000080)     //  syndrome : 0x09d4
                                | ({32{i_sel[144]}} & 32'h00000080)     //  syndrome : 0x09d7
                                | ({32{i_sel[143]}} & 32'h00000060)     //  syndrome : 0x0c03
                                | ({32{i_sel[142]}} & 32'h00000050)     //  syndrome : 0x1f3b
                                | ({32{i_sel[141]}} & 32'h00000048)     //  syndrome : 0x16a7
                                | ({32{i_sel[140]}} & 32'h00000044)     //  syndrome : 0x1269
                                | ({32{i_sel[139]}} & 32'h00000042)     //  syndrome : 0x0536
                                | ({32{i_sel[138]}} & 32'h00000041)     //  syndrome : 0x1ba0
                                | ({32{i_sel[137]}} & 32'h00000040)     //  syndrome : 0x01d3
                                | ({32{i_sel[136]}} & 32'h00000040)     //  syndrome : 0x19d3
                                | ({32{i_sel[135]}} & 32'h00000040)     //  syndrome : 0x15d3
                                | ({32{i_sel[134]}} & 32'h00000040)     //  syndrome : 0x13d3
                                | ({32{i_sel[133]}} & 32'h00000040)     //  syndrome : 0x10d3
                                | ({32{i_sel[132]}} & 32'h00000040)     //  syndrome : 0x1153
                                | ({32{i_sel[131]}} & 32'h00000040)     //  syndrome : 0x1193
                                | ({32{i_sel[130]}} & 32'h00000040)     //  syndrome : 0x11f3
                                | ({32{i_sel[129]}} & 32'h00000040)     //  syndrome : 0x11c3
                                | ({32{i_sel[128]}} & 32'h00000040)     //  syndrome : 0x11db
                                | ({32{i_sel[127]}} & 32'h00000040)     //  syndrome : 0x11d7
                                | ({32{i_sel[126]}} & 32'h00000040)     //  syndrome : 0x11d1
                                | ({32{i_sel[125]}} & 32'h00000040)     //  syndrome : 0x11d2
                                | ({32{i_sel[124]}} & 32'h00000030)     //  syndrome : 0x1338
                                | ({32{i_sel[123]}} & 32'h00000028)     //  syndrome : 0x1aa4
                                | ({32{i_sel[122]}} & 32'h00000024)     //  syndrome : 0x1e6a
                                | ({32{i_sel[121]}} & 32'h00000022)     //  syndrome : 0x0935
                                | ({32{i_sel[120]}} & 32'h00000021)     //  syndrome : 0x17a3
                                | ({32{i_sel[119]}} & 32'h00000020)     //  syndrome : 0x0dd0
                                | ({32{i_sel[118]}} & 32'h00000020)     //  syndrome : 0x15d0
                                | ({32{i_sel[117]}} & 32'h00000020)     //  syndrome : 0x19d0
                                | ({32{i_sel[116]}} & 32'h00000020)     //  syndrome : 0x1fd0
                                | ({32{i_sel[115]}} & 32'h00000020)     //  syndrome : 0x1cd0
                                | ({32{i_sel[114]}} & 32'h00000020)     //  syndrome : 0x1d50
                                | ({32{i_sel[113]}} & 32'h00000020)     //  syndrome : 0x1d90
                                | ({32{i_sel[112]}} & 32'h00000020)     //  syndrome : 0x1df0
                                | ({32{i_sel[111]}} & 32'h00000020)     //  syndrome : 0x1dc0
                                | ({32{i_sel[110]}} & 32'h00000020)     //  syndrome : 0x1dd8
                                | ({32{i_sel[109]}} & 32'h00000020)     //  syndrome : 0x1dd4
                                | ({32{i_sel[108]}} & 32'h00000020)     //  syndrome : 0x1dd2
                                | ({32{i_sel[107]}} & 32'h00000020)     //  syndrome : 0x1dd1
                                | ({32{i_sel[106]}} & 32'h00000018)     //  syndrome : 0x099c
                                | ({32{i_sel[105]}} & 32'h00000014)     //  syndrome : 0x0d52
                                | ({32{i_sel[104]}} & 32'h00000012)     //  syndrome : 0x1a0d
                                | ({32{i_sel[103]}} & 32'h00000011)     //  syndrome : 0x049b
                                | ({32{i_sel[102]}} & 32'h00000010)     //  syndrome : 0x1ee8
                                | ({32{i_sel[101]}} & 32'h00000010)     //  syndrome : 0x06e8
                                | ({32{i_sel[100]}} & 32'h00000010)     //  syndrome : 0x0ae8
                                | ({32{i_sel[99 ]}} & 32'h00000010)     //  syndrome : 0x0ce8
                                | ({32{i_sel[98 ]}} & 32'h00000010)     //  syndrome : 0x0fe8
                                | ({32{i_sel[97 ]}} & 32'h00000010)     //  syndrome : 0x0e68
                                | ({32{i_sel[96 ]}} & 32'h00000010)     //  syndrome : 0x0ea8
                                | ({32{i_sel[95 ]}} & 32'h00000010)     //  syndrome : 0x0ec8
                                | ({32{i_sel[94 ]}} & 32'h00000010)     //  syndrome : 0x0ef8
                                | ({32{i_sel[93 ]}} & 32'h00000010)     //  syndrome : 0x0ee0
                                | ({32{i_sel[92 ]}} & 32'h00000010)     //  syndrome : 0x0eec
                                | ({32{i_sel[91 ]}} & 32'h00000010)     //  syndrome : 0x0eea
                                | ({32{i_sel[90 ]}} & 32'h00000010)     //  syndrome : 0x0ee9
                                | ({32{i_sel[89 ]}} & 32'h0000000c)     //  syndrome : 0x04ce
                                | ({32{i_sel[88 ]}} & 32'h0000000a)     //  syndrome : 0x1391
                                | ({32{i_sel[87 ]}} & 32'h00000009)     //  syndrome : 0x0d07
                                | ({32{i_sel[86 ]}} & 32'h00000008)     //  syndrome : 0x1774
                                | ({32{i_sel[85 ]}} & 32'h00000008)     //  syndrome : 0x0f74
                                | ({32{i_sel[84 ]}} & 32'h00000008)     //  syndrome : 0x0374
                                | ({32{i_sel[83 ]}} & 32'h00000008)     //  syndrome : 0x0574
                                | ({32{i_sel[82 ]}} & 32'h00000008)     //  syndrome : 0x0674
                                | ({32{i_sel[81 ]}} & 32'h00000008)     //  syndrome : 0x07f4
                                | ({32{i_sel[80 ]}} & 32'h00000008)     //  syndrome : 0x0734
                                | ({32{i_sel[79 ]}} & 32'h00000008)     //  syndrome : 0x0754
                                | ({32{i_sel[78 ]}} & 32'h00000008)     //  syndrome : 0x0764
                                | ({32{i_sel[77 ]}} & 32'h00000008)     //  syndrome : 0x077c
                                | ({32{i_sel[76 ]}} & 32'h00000008)     //  syndrome : 0x0770
                                | ({32{i_sel[75 ]}} & 32'h00000008)     //  syndrome : 0x0776
                                | ({32{i_sel[74 ]}} & 32'h00000008)     //  syndrome : 0x0775
                                | ({32{i_sel[73 ]}} & 32'h00000006)     //  syndrome : 0x175f
                                | ({32{i_sel[72 ]}} & 32'h00000005)     //  syndrome : 0x09c9
                                | ({32{i_sel[71 ]}} & 32'h00000004)     //  syndrome : 0x13ba
                                | ({32{i_sel[70 ]}} & 32'h00000004)     //  syndrome : 0x0bba
                                | ({32{i_sel[69 ]}} & 32'h00000004)     //  syndrome : 0x07ba
                                | ({32{i_sel[68 ]}} & 32'h00000004)     //  syndrome : 0x01ba
                                | ({32{i_sel[67 ]}} & 32'h00000004)     //  syndrome : 0x02ba
                                | ({32{i_sel[66 ]}} & 32'h00000004)     //  syndrome : 0x033a
                                | ({32{i_sel[65 ]}} & 32'h00000004)     //  syndrome : 0x03fa
                                | ({32{i_sel[64 ]}} & 32'h00000004)     //  syndrome : 0x039a
                                | ({32{i_sel[63 ]}} & 32'h00000004)     //  syndrome : 0x03aa
                                | ({32{i_sel[62 ]}} & 32'h00000004)     //  syndrome : 0x03b2
                                | ({32{i_sel[61 ]}} & 32'h00000004)     //  syndrome : 0x03be
                                | ({32{i_sel[60 ]}} & 32'h00000004)     //  syndrome : 0x03b8
                                | ({32{i_sel[59 ]}} & 32'h00000004)     //  syndrome : 0x03bb
                                | ({32{i_sel[58 ]}} & 32'h00000003)     //  syndrome : 0x1e96
                                | ({32{i_sel[57 ]}} & 32'h00000002)     //  syndrome : 0x04e5
                                | ({32{i_sel[56 ]}} & 32'h00000002)     //  syndrome : 0x1ce5
                                | ({32{i_sel[55 ]}} & 32'h00000002)     //  syndrome : 0x10e5
                                | ({32{i_sel[54 ]}} & 32'h00000002)     //  syndrome : 0x16e5
                                | ({32{i_sel[53 ]}} & 32'h00000002)     //  syndrome : 0x15e5
                                | ({32{i_sel[52 ]}} & 32'h00000002)     //  syndrome : 0x1465
                                | ({32{i_sel[51 ]}} & 32'h00000002)     //  syndrome : 0x14a5
                                | ({32{i_sel[50 ]}} & 32'h00000002)     //  syndrome : 0x14c5
                                | ({32{i_sel[49 ]}} & 32'h00000002)     //  syndrome : 0x14f5
                                | ({32{i_sel[48 ]}} & 32'h00000002)     //  syndrome : 0x14ed
                                | ({32{i_sel[47 ]}} & 32'h00000002)     //  syndrome : 0x14e1
                                | ({32{i_sel[46 ]}} & 32'h00000002)     //  syndrome : 0x14e7
                                | ({32{i_sel[45 ]}} & 32'h00000002)     //  syndrome : 0x14e4
                                | ({32{i_sel[44 ]}} & 32'h00000001)     //  syndrome : 0x1a73
                                | ({32{i_sel[43 ]}} & 32'h00000001)     //  syndrome : 0x0273
                                | ({32{i_sel[42 ]}} & 32'h00000001)     //  syndrome : 0x0e73
                                | ({32{i_sel[41 ]}} & 32'h00000001)     //  syndrome : 0x0873
                                | ({32{i_sel[40 ]}} & 32'h00000001)     //  syndrome : 0x0b73
                                | ({32{i_sel[39 ]}} & 32'h00000001)     //  syndrome : 0x0af3
                                | ({32{i_sel[38 ]}} & 32'h00000001)     //  syndrome : 0x0a33
                                | ({32{i_sel[37 ]}} & 32'h00000001)     //  syndrome : 0x0a53
                                | ({32{i_sel[36 ]}} & 32'h00000001)     //  syndrome : 0x0a63
                                | ({32{i_sel[35 ]}} & 32'h00000001)     //  syndrome : 0x0a7b
                                | ({32{i_sel[34 ]}} & 32'h00000001)     //  syndrome : 0x0a77
                                | ({32{i_sel[33 ]}} & 32'h00000001)     //  syndrome : 0x0a71
                                | ({32{i_sel[32 ]}} & 32'h00000001)     //  syndrome : 0x0a72
                                | ({32{i_sel[31 ]}} & 32'h80000000)     //  syndrome : 0x07cc
                                | ({32{i_sel[30 ]}} & 32'h40000000)     //  syndrome : 0x03e6
                                | ({32{i_sel[29 ]}} & 32'h20000000)     //  syndrome : 0x14cb
                                | ({32{i_sel[28 ]}} & 32'h10000000)     //  syndrome : 0x1f5c
                                | ({32{i_sel[27 ]}} & 32'h08000000)     //  syndrome : 0x0fae
                                | ({32{i_sel[26 ]}} & 32'h04000000)     //  syndrome : 0x12ef
                                | ({32{i_sel[25 ]}} & 32'h02000000)     //  syndrome : 0x1c4e
                                | ({32{i_sel[24 ]}} & 32'h01000000)     //  syndrome : 0x1b1f
                                | ({32{i_sel[23 ]}} & 32'h00800000)     //  syndrome : 0x18b6
                                | ({32{i_sel[22 ]}} & 32'h00400000)     //  syndrome : 0x1963
                                | ({32{i_sel[21 ]}} & 32'h00200000)     //  syndrome : 0x1988
                                | ({32{i_sel[20 ]}} & 32'h00100000)     //  syndrome : 0x0cc4
                                | ({32{i_sel[19 ]}} & 32'h00080000)     //  syndrome : 0x0662
                                | ({32{i_sel[18 ]}} & 32'h00040000)     //  syndrome : 0x1609
                                | ({32{i_sel[17 ]}} & 32'h00020000)     //  syndrome : 0x0b05
                                | ({32{i_sel[16 ]}} & 32'h00010000)     //  syndrome : 0x0583
                                | ({32{i_sel[15 ]}} & 32'h00008000)     //  syndrome : 0x17f8
                                | ({32{i_sel[14 ]}} & 32'h00004000)     //  syndrome : 0x0bfc
                                | ({32{i_sel[13 ]}} & 32'h00002000)     //  syndrome : 0x05fe
                                | ({32{i_sel[12 ]}} & 32'h00001000)     //  syndrome : 0x17c7
                                | ({32{i_sel[11 ]}} & 32'h00000800)     //  syndrome : 0x1eda
                                | ({32{i_sel[10 ]}} & 32'h00000400)     //  syndrome : 0x1a55
                                | ({32{i_sel[9  ]}} & 32'h00000200)     //  syndrome : 0x0d2b
                                | ({32{i_sel[8  ]}} & 32'h00000100)     //  syndrome : 0x13ac
                                | ({32{i_sel[7  ]}} & 32'h00000080)     //  syndrome : 0x09d6
                                | ({32{i_sel[6  ]}} & 32'h00000040)     //  syndrome : 0x11d3
                                | ({32{i_sel[5  ]}} & 32'h00000020)     //  syndrome : 0x1dd0
                                | ({32{i_sel[4  ]}} & 32'h00000010)     //  syndrome : 0x0ee8
                                | ({32{i_sel[3  ]}} & 32'h00000008)     //  syndrome : 0x0774
                                | ({32{i_sel[2  ]}} & 32'h00000004)     //  syndrome : 0x03ba
                                | ({32{i_sel[1  ]}} & 32'h00000002)     //  syndrome : 0x14e5
                                | ({32{i_sel[0  ]}} & 32'h00000001);    //  syndrome : 0x0a73
endfunction
